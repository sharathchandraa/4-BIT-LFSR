magic
tech scmos
timestamp 1398581887
<< nwell >>
rect -1258 -15 -1230 10
rect -1190 -12 -1137 13
rect -1093 -12 -1040 13
rect -1007 -12 -954 13
rect -933 -12 -880 13
rect -779 -12 -726 13
rect -683 -12 -630 13
rect -601 -12 -548 13
rect -519 -12 -466 13
rect -1188 -93 -1160 -68
rect -777 -89 -749 -64
rect -1250 -195 -1222 -170
rect -1182 -192 -1129 -167
rect -1085 -192 -1032 -167
rect -999 -192 -946 -167
rect -925 -192 -872 -167
rect -771 -192 -718 -167
rect -675 -192 -622 -167
rect -593 -192 -540 -167
rect -511 -192 -458 -167
rect -1180 -273 -1152 -248
rect -769 -269 -741 -244
rect -1253 -371 -1225 -346
rect -1185 -368 -1132 -343
rect -1088 -368 -1035 -343
rect -1002 -368 -949 -343
rect -928 -368 -875 -343
rect -774 -368 -721 -343
rect -678 -368 -625 -343
rect -596 -368 -543 -343
rect -514 -368 -461 -343
rect -1183 -449 -1155 -424
rect -772 -445 -744 -420
rect -1245 -545 -1217 -520
rect -1177 -542 -1124 -517
rect -1080 -542 -1027 -517
rect -994 -542 -941 -517
rect -920 -542 -867 -517
rect -766 -542 -713 -517
rect -670 -542 -617 -517
rect -588 -542 -535 -517
rect -506 -542 -453 -517
rect -1175 -623 -1147 -598
rect -764 -619 -736 -594
<< polysilicon >>
rect -1179 2 -1177 4
rect -1151 2 -1149 4
rect -1082 2 -1080 4
rect -1054 2 -1052 4
rect -996 2 -994 4
rect -968 2 -966 4
rect -922 2 -920 4
rect -894 2 -892 4
rect -768 2 -766 4
rect -740 2 -738 4
rect -672 2 -670 4
rect -644 2 -642 4
rect -590 2 -588 4
rect -562 2 -560 4
rect -508 2 -506 4
rect -480 2 -478 4
rect -1245 0 -1243 2
rect -1245 -19 -1243 -8
rect -1248 -21 -1243 -19
rect -1245 -29 -1243 -21
rect -1179 -27 -1177 -6
rect -1151 -27 -1149 -6
rect -1082 -27 -1080 -6
rect -1054 -27 -1052 -6
rect -996 -27 -994 -6
rect -968 -27 -966 -6
rect -922 -27 -920 -6
rect -894 -27 -892 -6
rect -768 -27 -766 -6
rect -740 -27 -738 -6
rect -672 -27 -670 -6
rect -644 -27 -642 -6
rect -590 -27 -588 -6
rect -562 -27 -560 -6
rect -508 -27 -506 -6
rect -480 -27 -478 -6
rect -1179 -33 -1177 -31
rect -1151 -33 -1149 -31
rect -1082 -33 -1080 -31
rect -1054 -33 -1052 -31
rect -996 -33 -994 -31
rect -968 -33 -966 -31
rect -922 -33 -920 -31
rect -894 -33 -892 -31
rect -768 -33 -766 -31
rect -740 -33 -738 -31
rect -672 -33 -670 -31
rect -644 -33 -642 -31
rect -590 -33 -588 -31
rect -562 -33 -560 -31
rect -508 -33 -506 -31
rect -480 -33 -478 -31
rect -1245 -35 -1243 -33
rect -764 -74 -762 -72
rect -1175 -78 -1173 -76
rect -1175 -97 -1173 -86
rect -764 -93 -762 -82
rect -767 -95 -762 -93
rect -1178 -99 -1173 -97
rect -1175 -107 -1173 -99
rect -764 -103 -762 -95
rect -764 -109 -762 -107
rect -1175 -113 -1173 -111
rect -1171 -178 -1169 -176
rect -1143 -178 -1141 -176
rect -1074 -178 -1072 -176
rect -1046 -178 -1044 -176
rect -988 -178 -986 -176
rect -960 -178 -958 -176
rect -914 -178 -912 -176
rect -886 -178 -884 -176
rect -760 -178 -758 -176
rect -732 -178 -730 -176
rect -664 -178 -662 -176
rect -636 -178 -634 -176
rect -582 -178 -580 -176
rect -554 -178 -552 -176
rect -500 -178 -498 -176
rect -472 -178 -470 -176
rect -1237 -180 -1235 -178
rect -1237 -199 -1235 -188
rect -1240 -201 -1235 -199
rect -1237 -209 -1235 -201
rect -1171 -207 -1169 -186
rect -1143 -207 -1141 -186
rect -1074 -207 -1072 -186
rect -1046 -207 -1044 -186
rect -988 -207 -986 -186
rect -960 -207 -958 -186
rect -914 -207 -912 -186
rect -886 -207 -884 -186
rect -760 -207 -758 -186
rect -732 -207 -730 -186
rect -664 -207 -662 -186
rect -636 -207 -634 -186
rect -582 -207 -580 -186
rect -554 -207 -552 -186
rect -500 -207 -498 -186
rect -472 -207 -470 -186
rect -1171 -213 -1169 -211
rect -1143 -213 -1141 -211
rect -1074 -213 -1072 -211
rect -1046 -213 -1044 -211
rect -988 -213 -986 -211
rect -960 -213 -958 -211
rect -914 -213 -912 -211
rect -886 -213 -884 -211
rect -760 -213 -758 -211
rect -732 -213 -730 -211
rect -664 -213 -662 -211
rect -636 -213 -634 -211
rect -582 -213 -580 -211
rect -554 -213 -552 -211
rect -500 -213 -498 -211
rect -472 -213 -470 -211
rect -1237 -215 -1235 -213
rect -756 -254 -754 -252
rect -1167 -258 -1165 -256
rect -1167 -277 -1165 -266
rect -756 -273 -754 -262
rect -759 -275 -754 -273
rect -1170 -279 -1165 -277
rect -1167 -287 -1165 -279
rect -756 -283 -754 -275
rect -756 -289 -754 -287
rect -1167 -293 -1165 -291
rect -1174 -354 -1172 -352
rect -1146 -354 -1144 -352
rect -1077 -354 -1075 -352
rect -1049 -354 -1047 -352
rect -991 -354 -989 -352
rect -963 -354 -961 -352
rect -917 -354 -915 -352
rect -889 -354 -887 -352
rect -763 -354 -761 -352
rect -735 -354 -733 -352
rect -667 -354 -665 -352
rect -639 -354 -637 -352
rect -585 -354 -583 -352
rect -557 -354 -555 -352
rect -503 -354 -501 -352
rect -475 -354 -473 -352
rect -1240 -356 -1238 -354
rect -1240 -375 -1238 -364
rect -1243 -377 -1238 -375
rect -1240 -385 -1238 -377
rect -1174 -383 -1172 -362
rect -1146 -383 -1144 -362
rect -1077 -383 -1075 -362
rect -1049 -383 -1047 -362
rect -991 -383 -989 -362
rect -963 -383 -961 -362
rect -917 -383 -915 -362
rect -889 -383 -887 -362
rect -763 -383 -761 -362
rect -735 -383 -733 -362
rect -667 -383 -665 -362
rect -639 -383 -637 -362
rect -585 -383 -583 -362
rect -557 -383 -555 -362
rect -503 -383 -501 -362
rect -475 -383 -473 -362
rect -1174 -389 -1172 -387
rect -1146 -389 -1144 -387
rect -1077 -389 -1075 -387
rect -1049 -389 -1047 -387
rect -991 -389 -989 -387
rect -963 -389 -961 -387
rect -917 -389 -915 -387
rect -889 -389 -887 -387
rect -763 -389 -761 -387
rect -735 -389 -733 -387
rect -667 -389 -665 -387
rect -639 -389 -637 -387
rect -585 -389 -583 -387
rect -557 -389 -555 -387
rect -503 -389 -501 -387
rect -475 -389 -473 -387
rect -1240 -391 -1238 -389
rect -759 -430 -757 -428
rect -1170 -434 -1168 -432
rect -1170 -453 -1168 -442
rect -759 -449 -757 -438
rect -762 -451 -757 -449
rect -1173 -455 -1168 -453
rect -1170 -463 -1168 -455
rect -759 -459 -757 -451
rect -759 -465 -757 -463
rect -1170 -469 -1168 -467
rect -1166 -528 -1164 -526
rect -1138 -528 -1136 -526
rect -1069 -528 -1067 -526
rect -1041 -528 -1039 -526
rect -983 -528 -981 -526
rect -955 -528 -953 -526
rect -909 -528 -907 -526
rect -881 -528 -879 -526
rect -755 -528 -753 -526
rect -727 -528 -725 -526
rect -659 -528 -657 -526
rect -631 -528 -629 -526
rect -577 -528 -575 -526
rect -549 -528 -547 -526
rect -495 -528 -493 -526
rect -467 -528 -465 -526
rect -1232 -530 -1230 -528
rect -1232 -549 -1230 -538
rect -1235 -551 -1230 -549
rect -1232 -559 -1230 -551
rect -1166 -557 -1164 -536
rect -1138 -557 -1136 -536
rect -1069 -557 -1067 -536
rect -1041 -557 -1039 -536
rect -983 -557 -981 -536
rect -955 -557 -953 -536
rect -909 -557 -907 -536
rect -881 -557 -879 -536
rect -755 -557 -753 -536
rect -727 -557 -725 -536
rect -659 -557 -657 -536
rect -631 -557 -629 -536
rect -577 -557 -575 -536
rect -549 -557 -547 -536
rect -495 -557 -493 -536
rect -467 -557 -465 -536
rect -1166 -563 -1164 -561
rect -1138 -563 -1136 -561
rect -1069 -563 -1067 -561
rect -1041 -563 -1039 -561
rect -983 -563 -981 -561
rect -955 -563 -953 -561
rect -909 -563 -907 -561
rect -881 -563 -879 -561
rect -755 -563 -753 -561
rect -727 -563 -725 -561
rect -659 -563 -657 -561
rect -631 -563 -629 -561
rect -577 -563 -575 -561
rect -549 -563 -547 -561
rect -495 -563 -493 -561
rect -467 -563 -465 -561
rect -1232 -565 -1230 -563
rect -751 -604 -749 -602
rect -1162 -608 -1160 -606
rect -1162 -627 -1160 -616
rect -751 -623 -749 -612
rect -754 -625 -749 -623
rect -1165 -629 -1160 -627
rect -1162 -637 -1160 -629
rect -751 -633 -749 -625
rect -751 -639 -749 -637
rect -1162 -643 -1160 -641
<< ndiffusion >>
rect -1248 -33 -1245 -29
rect -1243 -33 -1240 -29
rect -1182 -31 -1179 -27
rect -1177 -31 -1174 -27
rect -1154 -31 -1151 -27
rect -1149 -31 -1146 -27
rect -1085 -31 -1082 -27
rect -1080 -31 -1077 -27
rect -1057 -31 -1054 -27
rect -1052 -31 -1049 -27
rect -999 -31 -996 -27
rect -994 -31 -991 -27
rect -971 -31 -968 -27
rect -966 -31 -963 -27
rect -925 -31 -922 -27
rect -920 -31 -917 -27
rect -897 -31 -894 -27
rect -892 -31 -889 -27
rect -771 -31 -768 -27
rect -766 -31 -763 -27
rect -743 -31 -740 -27
rect -738 -31 -735 -27
rect -675 -31 -672 -27
rect -670 -31 -667 -27
rect -647 -31 -644 -27
rect -642 -31 -639 -27
rect -593 -31 -590 -27
rect -588 -31 -585 -27
rect -565 -31 -562 -27
rect -560 -31 -557 -27
rect -511 -31 -508 -27
rect -506 -31 -503 -27
rect -483 -31 -480 -27
rect -478 -31 -475 -27
rect -1178 -111 -1175 -107
rect -1173 -111 -1170 -107
rect -767 -107 -764 -103
rect -762 -107 -759 -103
rect -1240 -213 -1237 -209
rect -1235 -213 -1232 -209
rect -1174 -211 -1171 -207
rect -1169 -211 -1166 -207
rect -1146 -211 -1143 -207
rect -1141 -211 -1138 -207
rect -1077 -211 -1074 -207
rect -1072 -211 -1069 -207
rect -1049 -211 -1046 -207
rect -1044 -211 -1041 -207
rect -991 -211 -988 -207
rect -986 -211 -983 -207
rect -963 -211 -960 -207
rect -958 -211 -955 -207
rect -917 -211 -914 -207
rect -912 -211 -909 -207
rect -889 -211 -886 -207
rect -884 -211 -881 -207
rect -763 -211 -760 -207
rect -758 -211 -755 -207
rect -735 -211 -732 -207
rect -730 -211 -727 -207
rect -667 -211 -664 -207
rect -662 -211 -659 -207
rect -639 -211 -636 -207
rect -634 -211 -631 -207
rect -585 -211 -582 -207
rect -580 -211 -577 -207
rect -557 -211 -554 -207
rect -552 -211 -549 -207
rect -503 -211 -500 -207
rect -498 -211 -495 -207
rect -475 -211 -472 -207
rect -470 -211 -467 -207
rect -1170 -291 -1167 -287
rect -1165 -291 -1162 -287
rect -759 -287 -756 -283
rect -754 -287 -751 -283
rect -1243 -389 -1240 -385
rect -1238 -389 -1235 -385
rect -1177 -387 -1174 -383
rect -1172 -387 -1169 -383
rect -1149 -387 -1146 -383
rect -1144 -387 -1141 -383
rect -1080 -387 -1077 -383
rect -1075 -387 -1072 -383
rect -1052 -387 -1049 -383
rect -1047 -387 -1044 -383
rect -994 -387 -991 -383
rect -989 -387 -986 -383
rect -966 -387 -963 -383
rect -961 -387 -958 -383
rect -920 -387 -917 -383
rect -915 -387 -912 -383
rect -892 -387 -889 -383
rect -887 -387 -884 -383
rect -766 -387 -763 -383
rect -761 -387 -758 -383
rect -738 -387 -735 -383
rect -733 -387 -730 -383
rect -670 -387 -667 -383
rect -665 -387 -662 -383
rect -642 -387 -639 -383
rect -637 -387 -634 -383
rect -588 -387 -585 -383
rect -583 -387 -580 -383
rect -560 -387 -557 -383
rect -555 -387 -552 -383
rect -506 -387 -503 -383
rect -501 -387 -498 -383
rect -478 -387 -475 -383
rect -473 -387 -470 -383
rect -1173 -467 -1170 -463
rect -1168 -467 -1165 -463
rect -762 -463 -759 -459
rect -757 -463 -754 -459
rect -1235 -563 -1232 -559
rect -1230 -563 -1227 -559
rect -1169 -561 -1166 -557
rect -1164 -561 -1161 -557
rect -1141 -561 -1138 -557
rect -1136 -561 -1133 -557
rect -1072 -561 -1069 -557
rect -1067 -561 -1064 -557
rect -1044 -561 -1041 -557
rect -1039 -561 -1036 -557
rect -986 -561 -983 -557
rect -981 -561 -978 -557
rect -958 -561 -955 -557
rect -953 -561 -950 -557
rect -912 -561 -909 -557
rect -907 -561 -904 -557
rect -884 -561 -881 -557
rect -879 -561 -876 -557
rect -758 -561 -755 -557
rect -753 -561 -750 -557
rect -730 -561 -727 -557
rect -725 -561 -722 -557
rect -662 -561 -659 -557
rect -657 -561 -654 -557
rect -634 -561 -631 -557
rect -629 -561 -626 -557
rect -580 -561 -577 -557
rect -575 -561 -572 -557
rect -552 -561 -549 -557
rect -547 -561 -544 -557
rect -498 -561 -495 -557
rect -493 -561 -490 -557
rect -470 -561 -467 -557
rect -465 -561 -462 -557
rect -1165 -641 -1162 -637
rect -1160 -641 -1157 -637
rect -754 -637 -751 -633
rect -749 -637 -746 -633
<< pdiffusion >>
rect -1248 -8 -1245 0
rect -1243 -8 -1240 0
rect -1181 -6 -1179 2
rect -1177 -6 -1175 2
rect -1153 -6 -1151 2
rect -1149 -6 -1147 2
rect -1084 -6 -1082 2
rect -1080 -6 -1078 2
rect -1056 -6 -1054 2
rect -1052 -6 -1050 2
rect -998 -6 -996 2
rect -994 -6 -992 2
rect -970 -6 -968 2
rect -966 -6 -964 2
rect -924 -6 -922 2
rect -920 -6 -918 2
rect -896 -6 -894 2
rect -892 -6 -890 2
rect -770 -6 -768 2
rect -766 -6 -764 2
rect -742 -6 -740 2
rect -738 -6 -736 2
rect -674 -6 -672 2
rect -670 -6 -668 2
rect -646 -6 -644 2
rect -642 -6 -640 2
rect -592 -6 -590 2
rect -588 -6 -586 2
rect -564 -6 -562 2
rect -560 -6 -558 2
rect -510 -6 -508 2
rect -506 -6 -504 2
rect -482 -6 -480 2
rect -478 -6 -476 2
rect -1178 -86 -1175 -78
rect -1173 -86 -1170 -78
rect -767 -82 -764 -74
rect -762 -82 -759 -74
rect -1240 -188 -1237 -180
rect -1235 -188 -1232 -180
rect -1173 -186 -1171 -178
rect -1169 -186 -1167 -178
rect -1145 -186 -1143 -178
rect -1141 -186 -1139 -178
rect -1076 -186 -1074 -178
rect -1072 -186 -1070 -178
rect -1048 -186 -1046 -178
rect -1044 -186 -1042 -178
rect -990 -186 -988 -178
rect -986 -186 -984 -178
rect -962 -186 -960 -178
rect -958 -186 -956 -178
rect -916 -186 -914 -178
rect -912 -186 -910 -178
rect -888 -186 -886 -178
rect -884 -186 -882 -178
rect -762 -186 -760 -178
rect -758 -186 -756 -178
rect -734 -186 -732 -178
rect -730 -186 -728 -178
rect -666 -186 -664 -178
rect -662 -186 -660 -178
rect -638 -186 -636 -178
rect -634 -186 -632 -178
rect -584 -186 -582 -178
rect -580 -186 -578 -178
rect -556 -186 -554 -178
rect -552 -186 -550 -178
rect -502 -186 -500 -178
rect -498 -186 -496 -178
rect -474 -186 -472 -178
rect -470 -186 -468 -178
rect -1170 -266 -1167 -258
rect -1165 -266 -1162 -258
rect -759 -262 -756 -254
rect -754 -262 -751 -254
rect -1243 -364 -1240 -356
rect -1238 -364 -1235 -356
rect -1176 -362 -1174 -354
rect -1172 -362 -1170 -354
rect -1148 -362 -1146 -354
rect -1144 -362 -1142 -354
rect -1079 -362 -1077 -354
rect -1075 -362 -1073 -354
rect -1051 -362 -1049 -354
rect -1047 -362 -1045 -354
rect -993 -362 -991 -354
rect -989 -362 -987 -354
rect -965 -362 -963 -354
rect -961 -362 -959 -354
rect -919 -362 -917 -354
rect -915 -362 -913 -354
rect -891 -362 -889 -354
rect -887 -362 -885 -354
rect -765 -362 -763 -354
rect -761 -362 -759 -354
rect -737 -362 -735 -354
rect -733 -362 -731 -354
rect -669 -362 -667 -354
rect -665 -362 -663 -354
rect -641 -362 -639 -354
rect -637 -362 -635 -354
rect -587 -362 -585 -354
rect -583 -362 -581 -354
rect -559 -362 -557 -354
rect -555 -362 -553 -354
rect -505 -362 -503 -354
rect -501 -362 -499 -354
rect -477 -362 -475 -354
rect -473 -362 -471 -354
rect -1173 -442 -1170 -434
rect -1168 -442 -1165 -434
rect -762 -438 -759 -430
rect -757 -438 -754 -430
rect -1235 -538 -1232 -530
rect -1230 -538 -1227 -530
rect -1168 -536 -1166 -528
rect -1164 -536 -1162 -528
rect -1140 -536 -1138 -528
rect -1136 -536 -1134 -528
rect -1071 -536 -1069 -528
rect -1067 -536 -1065 -528
rect -1043 -536 -1041 -528
rect -1039 -536 -1037 -528
rect -985 -536 -983 -528
rect -981 -536 -979 -528
rect -957 -536 -955 -528
rect -953 -536 -951 -528
rect -911 -536 -909 -528
rect -907 -536 -905 -528
rect -883 -536 -881 -528
rect -879 -536 -877 -528
rect -757 -536 -755 -528
rect -753 -536 -751 -528
rect -729 -536 -727 -528
rect -725 -536 -723 -528
rect -661 -536 -659 -528
rect -657 -536 -655 -528
rect -633 -536 -631 -528
rect -629 -536 -627 -528
rect -579 -536 -577 -528
rect -575 -536 -573 -528
rect -551 -536 -549 -528
rect -547 -536 -545 -528
rect -497 -536 -495 -528
rect -493 -536 -491 -528
rect -469 -536 -467 -528
rect -465 -536 -463 -528
rect -1165 -616 -1162 -608
rect -1160 -616 -1157 -608
rect -754 -612 -751 -604
rect -749 -612 -746 -604
<< metal1 >>
rect -1362 20 -492 23
rect -1362 -157 -1359 20
rect -1300 8 -1296 20
rect -1237 9 -1233 20
rect -1248 5 -1237 9
rect -1252 0 -1248 5
rect -1240 -18 -1236 -8
rect -1221 -18 -1217 11
rect -1167 10 -1163 20
rect -1070 10 -1066 20
rect -984 10 -980 20
rect -910 10 -906 20
rect -1181 6 -1177 10
rect -1173 6 -1167 10
rect -1163 6 -1157 10
rect -1153 6 -1147 10
rect -1185 2 -1181 6
rect -1147 2 -1143 6
rect -1171 -6 -1157 2
rect -1084 6 -1080 10
rect -1076 6 -1070 10
rect -1066 6 -1060 10
rect -1056 6 -1050 10
rect -1088 2 -1084 6
rect -1050 2 -1046 6
rect -1074 -6 -1060 2
rect -998 6 -994 10
rect -990 6 -984 10
rect -980 6 -974 10
rect -970 6 -964 10
rect -1002 2 -998 6
rect -964 2 -960 6
rect -988 -6 -974 2
rect -924 6 -920 10
rect -916 6 -910 10
rect -906 6 -900 10
rect -896 6 -890 10
rect -928 2 -924 6
rect -890 2 -886 6
rect -833 8 -829 20
rect -756 10 -752 20
rect -660 10 -656 20
rect -578 10 -574 20
rect -496 10 -492 20
rect -770 6 -766 10
rect -762 6 -756 10
rect -752 6 -746 10
rect -742 6 -736 10
rect -914 -6 -900 2
rect -1265 -22 -1252 -18
rect -1240 -22 -1217 -18
rect -1201 -18 -1183 -14
rect -1240 -28 -1236 -22
rect -1252 -38 -1248 -33
rect -1201 -36 -1197 -18
rect -1166 -21 -1163 -6
rect -1125 -14 -1121 -10
rect -1145 -18 -1121 -14
rect -1100 -18 -1086 -14
rect -1069 -21 -1066 -6
rect -1028 -14 -1024 -10
rect -1048 -18 -1024 -14
rect -1017 -18 -1000 -14
rect -1017 -21 -1014 -18
rect -983 -21 -980 -6
rect -950 -14 -946 -10
rect -962 -18 -946 -14
rect -938 -18 -926 -14
rect -938 -21 -935 -18
rect -909 -21 -906 -6
rect -888 -18 -878 -14
rect -1186 -24 -1118 -21
rect -1186 -27 -1182 -24
rect -1089 -24 -1014 -21
rect -1003 -24 -935 -21
rect -929 -24 -878 -21
rect -1089 -27 -1085 -24
rect -1003 -27 -999 -24
rect -929 -27 -925 -24
rect -1170 -32 -1158 -27
rect -1073 -32 -1061 -27
rect -987 -32 -975 -27
rect -913 -32 -901 -27
rect -881 -28 -878 -24
rect -869 -28 -864 -1
rect -774 2 -770 6
rect -736 2 -732 6
rect -760 -6 -746 2
rect -674 6 -670 10
rect -666 6 -660 10
rect -656 6 -650 10
rect -646 6 -640 10
rect -678 2 -674 6
rect -640 2 -636 6
rect -664 -6 -650 2
rect -592 6 -588 10
rect -584 6 -578 10
rect -574 6 -568 10
rect -564 6 -558 10
rect -596 2 -592 6
rect -558 2 -554 6
rect -582 -6 -568 2
rect -510 6 -506 10
rect -502 6 -496 10
rect -492 6 -486 10
rect -482 6 -476 10
rect -514 2 -510 6
rect -476 2 -472 6
rect -500 -6 -486 2
rect -790 -18 -772 -14
rect -790 -28 -786 -18
rect -755 -21 -752 -6
rect -714 -14 -710 -10
rect -734 -18 -710 -14
rect -690 -18 -676 -14
rect -659 -21 -656 -6
rect -618 -14 -614 -10
rect -638 -18 -614 -14
rect -605 -18 -594 -14
rect -605 -21 -602 -18
rect -577 -21 -574 -6
rect -536 -14 -532 -10
rect -556 -18 -532 -14
rect -525 -18 -512 -14
rect -525 -21 -522 -18
rect -495 -21 -492 -6
rect -474 -18 -464 -14
rect -881 -31 -786 -28
rect -1146 -37 -1142 -32
rect -1252 -45 -1248 -42
rect -1146 -45 -1142 -41
rect -1049 -37 -1045 -32
rect -1049 -45 -1045 -41
rect -963 -37 -959 -32
rect -963 -45 -959 -41
rect -889 -37 -885 -32
rect -790 -36 -786 -31
rect -775 -24 -706 -21
rect -775 -27 -771 -24
rect -679 -24 -602 -21
rect -597 -24 -522 -21
rect -515 -24 -464 -21
rect -679 -27 -675 -24
rect -597 -27 -593 -24
rect -515 -27 -511 -24
rect -759 -32 -747 -27
rect -663 -32 -651 -27
rect -581 -32 -569 -27
rect -499 -32 -487 -27
rect -467 -28 -464 -24
rect -455 -27 -450 -1
rect -455 -28 -363 -27
rect -467 -31 -363 -28
rect -735 -37 -731 -32
rect -889 -45 -885 -41
rect -735 -45 -731 -41
rect -639 -37 -635 -32
rect -639 -45 -635 -41
rect -557 -37 -553 -32
rect -557 -45 -553 -41
rect -475 -37 -471 -32
rect -475 -45 -471 -41
rect -1351 -48 -471 -45
rect -1351 -120 -1347 -48
rect -1319 -59 -1287 -54
rect -1319 -146 -1316 -59
rect -1234 -123 -1230 -48
rect -1148 -55 -1104 -51
rect -1213 -96 -1209 -65
rect -1196 -73 -1182 -69
rect -1178 -73 -1167 -69
rect -1182 -78 -1178 -73
rect -1170 -96 -1166 -86
rect -1148 -96 -1145 -55
rect -1213 -100 -1182 -96
rect -1170 -100 -1145 -96
rect -1170 -106 -1166 -100
rect -1182 -116 -1178 -111
rect -1182 -123 -1178 -120
rect -823 -119 -819 -48
rect -731 -55 -694 -51
rect -802 -92 -798 -59
rect -785 -69 -771 -65
rect -767 -69 -756 -65
rect -771 -74 -767 -69
rect -759 -92 -755 -82
rect -731 -92 -727 -55
rect -802 -96 -771 -92
rect -759 -96 -727 -92
rect -759 -102 -755 -96
rect -771 -112 -767 -107
rect -771 -119 -767 -116
rect -823 -122 -767 -119
rect -1234 -126 -1178 -123
rect -1319 -149 -423 -146
rect -1362 -160 -484 -157
rect -1362 -333 -1359 -160
rect -1292 -172 -1288 -160
rect -1229 -171 -1225 -160
rect -1240 -175 -1229 -171
rect -1244 -180 -1240 -175
rect -1232 -198 -1228 -188
rect -1213 -198 -1209 -169
rect -1159 -170 -1155 -160
rect -1062 -170 -1058 -160
rect -976 -170 -972 -160
rect -902 -170 -898 -160
rect -1173 -174 -1169 -170
rect -1165 -174 -1159 -170
rect -1155 -174 -1149 -170
rect -1145 -174 -1139 -170
rect -1177 -178 -1173 -174
rect -1139 -178 -1135 -174
rect -1163 -186 -1149 -178
rect -1076 -174 -1072 -170
rect -1068 -174 -1062 -170
rect -1058 -174 -1052 -170
rect -1048 -174 -1042 -170
rect -1080 -178 -1076 -174
rect -1042 -178 -1038 -174
rect -1066 -186 -1052 -178
rect -990 -174 -986 -170
rect -982 -174 -976 -170
rect -972 -174 -966 -170
rect -962 -174 -956 -170
rect -994 -178 -990 -174
rect -956 -178 -952 -174
rect -980 -186 -966 -178
rect -916 -174 -912 -170
rect -908 -174 -902 -170
rect -898 -174 -892 -170
rect -888 -174 -882 -170
rect -920 -178 -916 -174
rect -882 -178 -878 -174
rect -825 -172 -821 -160
rect -748 -170 -744 -160
rect -652 -170 -648 -160
rect -570 -170 -566 -160
rect -488 -170 -484 -160
rect -762 -174 -758 -170
rect -754 -174 -748 -170
rect -744 -174 -738 -170
rect -734 -174 -728 -170
rect -906 -186 -892 -178
rect -1257 -202 -1244 -198
rect -1232 -202 -1209 -198
rect -1193 -198 -1175 -194
rect -1232 -208 -1228 -202
rect -1244 -218 -1240 -213
rect -1193 -216 -1189 -198
rect -1158 -201 -1155 -186
rect -1117 -194 -1113 -190
rect -1137 -198 -1113 -194
rect -1092 -198 -1078 -194
rect -1061 -201 -1058 -186
rect -1020 -194 -1016 -190
rect -1040 -198 -1016 -194
rect -1009 -198 -992 -194
rect -1009 -201 -1006 -198
rect -975 -201 -972 -186
rect -942 -194 -938 -190
rect -954 -198 -938 -194
rect -930 -198 -918 -194
rect -930 -201 -927 -198
rect -901 -201 -898 -186
rect -880 -198 -870 -194
rect -1178 -204 -1110 -201
rect -1178 -207 -1174 -204
rect -1081 -204 -1006 -201
rect -995 -204 -927 -201
rect -921 -204 -870 -201
rect -1081 -207 -1077 -204
rect -995 -207 -991 -204
rect -921 -207 -917 -204
rect -1162 -212 -1150 -207
rect -1065 -212 -1053 -207
rect -979 -212 -967 -207
rect -905 -212 -893 -207
rect -873 -208 -870 -204
rect -861 -208 -856 -181
rect -766 -178 -762 -174
rect -728 -178 -724 -174
rect -752 -186 -738 -178
rect -666 -174 -662 -170
rect -658 -174 -652 -170
rect -648 -174 -642 -170
rect -638 -174 -632 -170
rect -670 -178 -666 -174
rect -632 -178 -628 -174
rect -656 -186 -642 -178
rect -584 -174 -580 -170
rect -576 -174 -570 -170
rect -566 -174 -560 -170
rect -556 -174 -550 -170
rect -588 -178 -584 -174
rect -550 -178 -546 -174
rect -574 -186 -560 -178
rect -502 -174 -498 -170
rect -494 -174 -488 -170
rect -484 -174 -478 -170
rect -474 -174 -468 -170
rect -506 -178 -502 -174
rect -468 -178 -464 -174
rect -492 -186 -478 -178
rect -782 -198 -764 -194
rect -782 -208 -778 -198
rect -747 -201 -744 -186
rect -706 -194 -702 -190
rect -726 -198 -702 -194
rect -682 -198 -668 -194
rect -651 -201 -648 -186
rect -610 -194 -606 -190
rect -630 -198 -606 -194
rect -597 -198 -586 -194
rect -597 -201 -594 -198
rect -569 -201 -566 -186
rect -528 -194 -524 -190
rect -548 -198 -524 -194
rect -517 -198 -504 -194
rect -517 -201 -514 -198
rect -487 -201 -484 -186
rect -466 -198 -456 -194
rect -873 -211 -778 -208
rect -1138 -217 -1134 -212
rect -1244 -225 -1240 -222
rect -1138 -225 -1134 -221
rect -1041 -217 -1037 -212
rect -1041 -225 -1037 -221
rect -955 -217 -951 -212
rect -955 -225 -951 -221
rect -881 -217 -877 -212
rect -782 -216 -778 -211
rect -767 -204 -698 -201
rect -767 -207 -763 -204
rect -671 -204 -594 -201
rect -589 -204 -514 -201
rect -507 -204 -456 -201
rect -671 -207 -667 -204
rect -589 -207 -585 -204
rect -507 -207 -503 -204
rect -751 -212 -739 -207
rect -655 -212 -643 -207
rect -573 -212 -561 -207
rect -491 -212 -479 -207
rect -459 -208 -456 -204
rect -447 -207 -442 -181
rect -426 -207 -423 -149
rect -447 -208 -423 -207
rect -459 -211 -423 -208
rect -727 -217 -723 -212
rect -881 -225 -877 -221
rect -727 -225 -723 -221
rect -631 -217 -627 -212
rect -631 -225 -627 -221
rect -549 -217 -545 -212
rect -549 -225 -545 -221
rect -467 -217 -463 -212
rect -467 -225 -463 -221
rect -1347 -228 -463 -225
rect -1316 -239 -1279 -234
rect -1316 -322 -1312 -239
rect -1226 -303 -1222 -228
rect -1140 -235 -1096 -231
rect -1205 -276 -1201 -245
rect -1188 -253 -1174 -249
rect -1170 -253 -1159 -249
rect -1174 -258 -1170 -253
rect -1162 -276 -1158 -266
rect -1140 -276 -1137 -235
rect -1205 -280 -1174 -276
rect -1162 -280 -1137 -276
rect -1162 -286 -1158 -280
rect -1174 -296 -1170 -291
rect -1174 -303 -1170 -300
rect -815 -299 -811 -228
rect -723 -235 -686 -231
rect -794 -272 -790 -239
rect -777 -249 -763 -245
rect -759 -249 -748 -245
rect -763 -254 -759 -249
rect -751 -272 -747 -262
rect -723 -272 -719 -235
rect -794 -276 -763 -272
rect -751 -276 -719 -272
rect -751 -282 -747 -276
rect -763 -292 -759 -287
rect -763 -299 -759 -296
rect -815 -302 -759 -299
rect -1226 -306 -1170 -303
rect -1316 -325 -425 -322
rect -1362 -336 -487 -333
rect -1362 -507 -1359 -336
rect -1295 -348 -1291 -336
rect -1232 -347 -1228 -336
rect -1243 -351 -1232 -347
rect -1247 -356 -1243 -351
rect -1235 -374 -1231 -364
rect -1216 -374 -1212 -345
rect -1162 -346 -1158 -336
rect -1065 -346 -1061 -336
rect -979 -346 -975 -336
rect -905 -346 -901 -336
rect -1176 -350 -1172 -346
rect -1168 -350 -1162 -346
rect -1158 -350 -1152 -346
rect -1148 -350 -1142 -346
rect -1180 -354 -1176 -350
rect -1142 -354 -1138 -350
rect -1166 -362 -1152 -354
rect -1079 -350 -1075 -346
rect -1071 -350 -1065 -346
rect -1061 -350 -1055 -346
rect -1051 -350 -1045 -346
rect -1083 -354 -1079 -350
rect -1045 -354 -1041 -350
rect -1069 -362 -1055 -354
rect -993 -350 -989 -346
rect -985 -350 -979 -346
rect -975 -350 -969 -346
rect -965 -350 -959 -346
rect -997 -354 -993 -350
rect -959 -354 -955 -350
rect -983 -362 -969 -354
rect -919 -350 -915 -346
rect -911 -350 -905 -346
rect -901 -350 -895 -346
rect -891 -350 -885 -346
rect -923 -354 -919 -350
rect -885 -354 -881 -350
rect -828 -348 -824 -336
rect -751 -346 -747 -336
rect -655 -346 -651 -336
rect -573 -346 -569 -336
rect -491 -346 -487 -336
rect -765 -350 -761 -346
rect -757 -350 -751 -346
rect -747 -350 -741 -346
rect -737 -350 -731 -346
rect -909 -362 -895 -354
rect -1260 -378 -1247 -374
rect -1235 -378 -1212 -374
rect -1196 -374 -1178 -370
rect -1235 -384 -1231 -378
rect -1247 -394 -1243 -389
rect -1196 -392 -1192 -374
rect -1161 -377 -1158 -362
rect -1120 -370 -1116 -366
rect -1140 -374 -1116 -370
rect -1095 -374 -1081 -370
rect -1064 -377 -1061 -362
rect -1023 -370 -1019 -366
rect -1043 -374 -1019 -370
rect -1012 -374 -995 -370
rect -1012 -377 -1009 -374
rect -978 -377 -975 -362
rect -945 -370 -941 -366
rect -957 -374 -941 -370
rect -933 -374 -921 -370
rect -933 -377 -930 -374
rect -904 -377 -901 -362
rect -883 -374 -873 -370
rect -1181 -380 -1113 -377
rect -1181 -383 -1177 -380
rect -1084 -380 -1009 -377
rect -998 -380 -930 -377
rect -924 -380 -873 -377
rect -1084 -383 -1080 -380
rect -998 -383 -994 -380
rect -924 -383 -920 -380
rect -1165 -388 -1153 -383
rect -1068 -388 -1056 -383
rect -982 -388 -970 -383
rect -908 -388 -896 -383
rect -876 -384 -873 -380
rect -864 -384 -859 -357
rect -769 -354 -765 -350
rect -731 -354 -727 -350
rect -755 -362 -741 -354
rect -669 -350 -665 -346
rect -661 -350 -655 -346
rect -651 -350 -645 -346
rect -641 -350 -635 -346
rect -673 -354 -669 -350
rect -635 -354 -631 -350
rect -659 -362 -645 -354
rect -587 -350 -583 -346
rect -579 -350 -573 -346
rect -569 -350 -563 -346
rect -559 -350 -553 -346
rect -591 -354 -587 -350
rect -553 -354 -549 -350
rect -577 -362 -563 -354
rect -505 -350 -501 -346
rect -497 -350 -491 -346
rect -487 -350 -481 -346
rect -477 -350 -471 -346
rect -509 -354 -505 -350
rect -471 -354 -467 -350
rect -495 -362 -481 -354
rect -785 -374 -767 -370
rect -785 -384 -781 -374
rect -750 -377 -747 -362
rect -709 -370 -705 -366
rect -729 -374 -705 -370
rect -685 -374 -671 -370
rect -654 -377 -651 -362
rect -613 -370 -609 -366
rect -633 -374 -609 -370
rect -600 -374 -589 -370
rect -600 -377 -597 -374
rect -572 -377 -569 -362
rect -531 -370 -527 -366
rect -551 -374 -527 -370
rect -520 -374 -507 -370
rect -520 -377 -517 -374
rect -490 -377 -487 -362
rect -469 -374 -459 -370
rect -876 -387 -781 -384
rect -1141 -393 -1137 -388
rect -1247 -401 -1243 -398
rect -1141 -401 -1137 -397
rect -1044 -393 -1040 -388
rect -1044 -401 -1040 -397
rect -958 -393 -954 -388
rect -958 -401 -954 -397
rect -884 -393 -880 -388
rect -785 -392 -781 -387
rect -770 -380 -701 -377
rect -770 -383 -766 -380
rect -674 -380 -597 -377
rect -592 -380 -517 -377
rect -510 -380 -459 -377
rect -674 -383 -670 -380
rect -592 -383 -588 -380
rect -510 -383 -506 -380
rect -754 -388 -742 -383
rect -658 -388 -646 -383
rect -576 -388 -564 -383
rect -494 -388 -482 -383
rect -462 -384 -459 -380
rect -450 -383 -445 -357
rect -428 -383 -425 -325
rect -450 -384 -425 -383
rect -462 -387 -425 -384
rect -730 -393 -726 -388
rect -884 -401 -880 -397
rect -730 -401 -726 -397
rect -634 -393 -630 -388
rect -634 -401 -630 -397
rect -552 -393 -548 -388
rect -552 -401 -548 -397
rect -470 -393 -466 -388
rect -470 -401 -466 -397
rect -1347 -404 -466 -401
rect -1315 -415 -1282 -410
rect -1315 -495 -1312 -415
rect -1229 -479 -1225 -404
rect -1143 -411 -1099 -407
rect -1208 -452 -1204 -421
rect -1191 -429 -1177 -425
rect -1173 -429 -1162 -425
rect -1177 -434 -1173 -429
rect -1165 -452 -1161 -442
rect -1143 -452 -1140 -411
rect -1208 -456 -1177 -452
rect -1165 -456 -1140 -452
rect -1165 -462 -1161 -456
rect -1177 -472 -1173 -467
rect -1177 -479 -1173 -476
rect -818 -475 -814 -404
rect -726 -411 -689 -407
rect -797 -448 -793 -415
rect -780 -425 -766 -421
rect -762 -425 -751 -421
rect -766 -430 -762 -425
rect -754 -448 -750 -438
rect -726 -448 -722 -411
rect -797 -452 -766 -448
rect -754 -452 -722 -448
rect -754 -458 -750 -452
rect -766 -468 -762 -463
rect -766 -475 -762 -472
rect -818 -478 -762 -475
rect -1229 -482 -1173 -479
rect -1315 -498 -417 -495
rect -1362 -510 -479 -507
rect -1362 -669 -1359 -510
rect -1287 -522 -1283 -510
rect -1224 -521 -1220 -510
rect -1235 -525 -1224 -521
rect -1239 -530 -1235 -525
rect -1227 -548 -1223 -538
rect -1208 -548 -1204 -519
rect -1154 -520 -1150 -510
rect -1057 -520 -1053 -510
rect -971 -520 -967 -510
rect -897 -520 -893 -510
rect -1168 -524 -1164 -520
rect -1160 -524 -1154 -520
rect -1150 -524 -1144 -520
rect -1140 -524 -1134 -520
rect -1172 -528 -1168 -524
rect -1134 -528 -1130 -524
rect -1158 -536 -1144 -528
rect -1071 -524 -1067 -520
rect -1063 -524 -1057 -520
rect -1053 -524 -1047 -520
rect -1043 -524 -1037 -520
rect -1075 -528 -1071 -524
rect -1037 -528 -1033 -524
rect -1061 -536 -1047 -528
rect -985 -524 -981 -520
rect -977 -524 -971 -520
rect -967 -524 -961 -520
rect -957 -524 -951 -520
rect -989 -528 -985 -524
rect -951 -528 -947 -524
rect -975 -536 -961 -528
rect -911 -524 -907 -520
rect -903 -524 -897 -520
rect -893 -524 -887 -520
rect -883 -524 -877 -520
rect -915 -528 -911 -524
rect -877 -528 -873 -524
rect -820 -522 -816 -510
rect -743 -520 -739 -510
rect -647 -520 -643 -510
rect -565 -520 -561 -510
rect -483 -520 -479 -510
rect -757 -524 -753 -520
rect -749 -524 -743 -520
rect -739 -524 -733 -520
rect -729 -524 -723 -520
rect -901 -536 -887 -528
rect -1252 -552 -1239 -548
rect -1227 -552 -1204 -548
rect -1188 -548 -1170 -544
rect -1227 -558 -1223 -552
rect -1239 -568 -1235 -563
rect -1188 -566 -1184 -548
rect -1153 -551 -1150 -536
rect -1112 -544 -1108 -540
rect -1132 -548 -1108 -544
rect -1087 -548 -1073 -544
rect -1056 -551 -1053 -536
rect -1015 -544 -1011 -540
rect -1035 -548 -1011 -544
rect -1004 -548 -987 -544
rect -1004 -551 -1001 -548
rect -970 -551 -967 -536
rect -937 -544 -933 -540
rect -949 -548 -933 -544
rect -925 -548 -913 -544
rect -925 -551 -922 -548
rect -896 -551 -893 -536
rect -875 -548 -865 -544
rect -1173 -554 -1105 -551
rect -1173 -557 -1169 -554
rect -1076 -554 -1001 -551
rect -990 -554 -922 -551
rect -916 -554 -865 -551
rect -1076 -557 -1072 -554
rect -990 -557 -986 -554
rect -916 -557 -912 -554
rect -1157 -562 -1145 -557
rect -1060 -562 -1048 -557
rect -974 -562 -962 -557
rect -900 -562 -888 -557
rect -868 -558 -865 -554
rect -856 -558 -851 -531
rect -761 -528 -757 -524
rect -723 -528 -719 -524
rect -747 -536 -733 -528
rect -661 -524 -657 -520
rect -653 -524 -647 -520
rect -643 -524 -637 -520
rect -633 -524 -627 -520
rect -665 -528 -661 -524
rect -627 -528 -623 -524
rect -651 -536 -637 -528
rect -579 -524 -575 -520
rect -571 -524 -565 -520
rect -561 -524 -555 -520
rect -551 -524 -545 -520
rect -583 -528 -579 -524
rect -545 -528 -541 -524
rect -569 -536 -555 -528
rect -497 -524 -493 -520
rect -489 -524 -483 -520
rect -479 -524 -473 -520
rect -469 -524 -463 -520
rect -501 -528 -497 -524
rect -463 -528 -459 -524
rect -487 -536 -473 -528
rect -777 -548 -759 -544
rect -777 -558 -773 -548
rect -742 -551 -739 -536
rect -701 -544 -697 -540
rect -721 -548 -697 -544
rect -677 -548 -663 -544
rect -646 -551 -643 -536
rect -605 -544 -601 -540
rect -625 -548 -601 -544
rect -592 -548 -581 -544
rect -592 -551 -589 -548
rect -564 -551 -561 -536
rect -523 -544 -519 -540
rect -543 -548 -519 -544
rect -512 -548 -499 -544
rect -512 -551 -509 -548
rect -482 -551 -479 -536
rect -461 -548 -451 -544
rect -868 -561 -773 -558
rect -1133 -567 -1129 -562
rect -1239 -575 -1235 -572
rect -1133 -575 -1129 -571
rect -1036 -567 -1032 -562
rect -1036 -575 -1032 -571
rect -950 -567 -946 -562
rect -950 -575 -946 -571
rect -876 -567 -872 -562
rect -777 -566 -773 -561
rect -762 -554 -693 -551
rect -762 -557 -758 -554
rect -666 -554 -589 -551
rect -584 -554 -509 -551
rect -502 -554 -451 -551
rect -666 -557 -662 -554
rect -584 -557 -580 -554
rect -502 -557 -498 -554
rect -746 -562 -734 -557
rect -650 -562 -638 -557
rect -568 -562 -556 -557
rect -486 -562 -474 -557
rect -454 -558 -451 -554
rect -442 -557 -437 -531
rect -420 -557 -417 -498
rect -442 -558 -417 -557
rect -454 -561 -417 -558
rect -722 -567 -718 -562
rect -876 -575 -872 -571
rect -722 -575 -718 -571
rect -626 -567 -622 -562
rect -626 -575 -622 -571
rect -544 -567 -540 -562
rect -544 -575 -540 -571
rect -462 -567 -458 -562
rect -462 -575 -458 -571
rect -1347 -578 -458 -575
rect -1304 -589 -1274 -584
rect -1221 -653 -1217 -578
rect -1135 -585 -1091 -581
rect -1200 -626 -1196 -595
rect -1183 -603 -1169 -599
rect -1165 -603 -1154 -599
rect -1169 -608 -1165 -603
rect -1157 -626 -1153 -616
rect -1135 -626 -1132 -585
rect -1200 -630 -1169 -626
rect -1157 -630 -1132 -626
rect -1157 -636 -1153 -630
rect -1169 -646 -1165 -641
rect -1169 -653 -1165 -650
rect -810 -649 -806 -578
rect -718 -585 -681 -581
rect -789 -622 -785 -589
rect -772 -599 -758 -595
rect -754 -599 -743 -595
rect -758 -604 -754 -599
rect -746 -622 -742 -612
rect -718 -622 -714 -585
rect -789 -626 -758 -622
rect -746 -626 -714 -622
rect -746 -632 -742 -626
rect -758 -642 -754 -637
rect -758 -649 -754 -646
rect -810 -652 -754 -649
rect -1221 -656 -1165 -653
rect -405 -727 -398 -31
<< metal2 >>
rect -1333 27 -614 30
rect -1351 -224 -1347 -124
rect -1351 -400 -1347 -228
rect -1351 -574 -1347 -404
rect -1351 -668 -1347 -578
rect -1333 -150 -1330 27
rect -1300 -69 -1296 4
rect -1270 -18 -1265 27
rect -1221 20 -1024 23
rect -1221 15 -1217 20
rect -1125 -6 -1121 20
rect -1028 -6 -1024 20
rect -950 20 -864 23
rect -950 -6 -946 20
rect -869 4 -864 20
rect -874 -18 -845 -14
rect -1213 -40 -1201 -36
rect -1213 -54 -1209 -40
rect -1282 -59 -1209 -54
rect -1213 -61 -1209 -59
rect -1118 -65 -1114 -25
rect -1104 -51 -1100 -18
rect -851 -65 -845 -18
rect -1118 -69 -845 -65
rect -833 -65 -829 4
rect -714 -6 -710 27
rect -618 -6 -614 27
rect -536 20 -450 23
rect -536 -6 -532 20
rect -455 4 -450 20
rect -460 -18 -436 -14
rect -802 -40 -790 -36
rect -802 -55 -798 -40
rect -706 -62 -702 -25
rect -694 -51 -690 -18
rect -442 -62 -436 -18
rect -833 -69 -789 -65
rect -706 -66 -436 -62
rect -1300 -73 -1200 -69
rect -1333 -153 -606 -150
rect -1333 -326 -1330 -153
rect -1292 -249 -1288 -176
rect -1262 -198 -1257 -153
rect -1213 -160 -1016 -157
rect -1213 -165 -1209 -160
rect -1117 -186 -1113 -160
rect -1020 -186 -1016 -160
rect -942 -160 -856 -157
rect -942 -186 -938 -160
rect -861 -176 -856 -160
rect -866 -198 -837 -194
rect -1205 -220 -1193 -216
rect -1205 -234 -1201 -220
rect -1274 -239 -1201 -234
rect -1205 -241 -1201 -239
rect -1110 -245 -1106 -205
rect -1096 -231 -1092 -198
rect -843 -245 -837 -198
rect -1110 -249 -837 -245
rect -825 -245 -821 -176
rect -706 -186 -702 -153
rect -610 -186 -606 -153
rect -528 -160 -442 -157
rect -528 -186 -524 -160
rect -447 -176 -442 -160
rect -452 -198 -428 -194
rect -794 -220 -782 -216
rect -794 -235 -790 -220
rect -698 -242 -694 -205
rect -686 -231 -682 -198
rect -434 -242 -428 -198
rect -419 -211 -362 -207
rect -825 -249 -781 -245
rect -698 -246 -428 -242
rect -1292 -253 -1192 -249
rect -1333 -329 -609 -326
rect -1333 -500 -1330 -329
rect -1295 -425 -1291 -352
rect -1265 -374 -1260 -329
rect -1216 -336 -1019 -333
rect -1216 -341 -1212 -336
rect -1120 -362 -1116 -336
rect -1023 -362 -1019 -336
rect -945 -336 -859 -333
rect -945 -362 -941 -336
rect -864 -352 -859 -336
rect -869 -374 -840 -370
rect -1208 -396 -1196 -392
rect -1208 -410 -1204 -396
rect -1277 -415 -1204 -410
rect -1208 -417 -1204 -415
rect -1113 -421 -1109 -381
rect -1099 -407 -1095 -374
rect -846 -421 -840 -374
rect -1113 -425 -840 -421
rect -828 -421 -824 -352
rect -709 -362 -705 -329
rect -613 -362 -609 -329
rect -531 -336 -445 -333
rect -531 -362 -527 -336
rect -450 -352 -445 -336
rect -455 -374 -431 -370
rect -797 -396 -785 -392
rect -797 -411 -793 -396
rect -701 -418 -697 -381
rect -689 -407 -685 -374
rect -437 -418 -431 -374
rect -421 -387 -360 -383
rect -828 -425 -784 -421
rect -701 -422 -431 -418
rect -1295 -429 -1195 -425
rect -1333 -503 -601 -500
rect -1333 -670 -1330 -503
rect -1287 -599 -1283 -526
rect -1257 -548 -1252 -503
rect -1208 -510 -1011 -507
rect -1208 -515 -1204 -510
rect -1112 -536 -1108 -510
rect -1015 -536 -1011 -510
rect -937 -510 -851 -507
rect -937 -536 -933 -510
rect -856 -526 -851 -510
rect -861 -548 -832 -544
rect -1200 -570 -1188 -566
rect -1200 -584 -1196 -570
rect -1269 -589 -1196 -584
rect -1200 -591 -1196 -589
rect -1105 -595 -1101 -555
rect -1091 -581 -1087 -548
rect -838 -595 -832 -548
rect -1105 -599 -832 -595
rect -820 -595 -816 -526
rect -701 -536 -697 -503
rect -605 -536 -601 -503
rect -523 -510 -437 -507
rect -523 -536 -519 -510
rect -442 -526 -437 -510
rect -447 -548 -423 -544
rect -789 -570 -777 -566
rect -789 -585 -785 -570
rect -693 -592 -689 -555
rect -681 -581 -677 -548
rect -429 -592 -423 -548
rect -413 -561 -371 -557
rect -820 -599 -776 -595
rect -693 -596 -423 -592
rect -1287 -603 -1187 -599
<< ntransistor >>
rect -1245 -33 -1243 -29
rect -1179 -31 -1177 -27
rect -1151 -31 -1149 -27
rect -1082 -31 -1080 -27
rect -1054 -31 -1052 -27
rect -996 -31 -994 -27
rect -968 -31 -966 -27
rect -922 -31 -920 -27
rect -894 -31 -892 -27
rect -768 -31 -766 -27
rect -740 -31 -738 -27
rect -672 -31 -670 -27
rect -644 -31 -642 -27
rect -590 -31 -588 -27
rect -562 -31 -560 -27
rect -508 -31 -506 -27
rect -480 -31 -478 -27
rect -1175 -111 -1173 -107
rect -764 -107 -762 -103
rect -1237 -213 -1235 -209
rect -1171 -211 -1169 -207
rect -1143 -211 -1141 -207
rect -1074 -211 -1072 -207
rect -1046 -211 -1044 -207
rect -988 -211 -986 -207
rect -960 -211 -958 -207
rect -914 -211 -912 -207
rect -886 -211 -884 -207
rect -760 -211 -758 -207
rect -732 -211 -730 -207
rect -664 -211 -662 -207
rect -636 -211 -634 -207
rect -582 -211 -580 -207
rect -554 -211 -552 -207
rect -500 -211 -498 -207
rect -472 -211 -470 -207
rect -1167 -291 -1165 -287
rect -756 -287 -754 -283
rect -1240 -389 -1238 -385
rect -1174 -387 -1172 -383
rect -1146 -387 -1144 -383
rect -1077 -387 -1075 -383
rect -1049 -387 -1047 -383
rect -991 -387 -989 -383
rect -963 -387 -961 -383
rect -917 -387 -915 -383
rect -889 -387 -887 -383
rect -763 -387 -761 -383
rect -735 -387 -733 -383
rect -667 -387 -665 -383
rect -639 -387 -637 -383
rect -585 -387 -583 -383
rect -557 -387 -555 -383
rect -503 -387 -501 -383
rect -475 -387 -473 -383
rect -1170 -467 -1168 -463
rect -759 -463 -757 -459
rect -1232 -563 -1230 -559
rect -1166 -561 -1164 -557
rect -1138 -561 -1136 -557
rect -1069 -561 -1067 -557
rect -1041 -561 -1039 -557
rect -983 -561 -981 -557
rect -955 -561 -953 -557
rect -909 -561 -907 -557
rect -881 -561 -879 -557
rect -755 -561 -753 -557
rect -727 -561 -725 -557
rect -659 -561 -657 -557
rect -631 -561 -629 -557
rect -577 -561 -575 -557
rect -549 -561 -547 -557
rect -495 -561 -493 -557
rect -467 -561 -465 -557
rect -1162 -641 -1160 -637
rect -751 -637 -749 -633
<< ptransistor >>
rect -1245 -8 -1243 0
rect -1179 -6 -1177 2
rect -1151 -6 -1149 2
rect -1082 -6 -1080 2
rect -1054 -6 -1052 2
rect -996 -6 -994 2
rect -968 -6 -966 2
rect -922 -6 -920 2
rect -894 -6 -892 2
rect -768 -6 -766 2
rect -740 -6 -738 2
rect -672 -6 -670 2
rect -644 -6 -642 2
rect -590 -6 -588 2
rect -562 -6 -560 2
rect -508 -6 -506 2
rect -480 -6 -478 2
rect -1175 -86 -1173 -78
rect -764 -82 -762 -74
rect -1237 -188 -1235 -180
rect -1171 -186 -1169 -178
rect -1143 -186 -1141 -178
rect -1074 -186 -1072 -178
rect -1046 -186 -1044 -178
rect -988 -186 -986 -178
rect -960 -186 -958 -178
rect -914 -186 -912 -178
rect -886 -186 -884 -178
rect -760 -186 -758 -178
rect -732 -186 -730 -178
rect -664 -186 -662 -178
rect -636 -186 -634 -178
rect -582 -186 -580 -178
rect -554 -186 -552 -178
rect -500 -186 -498 -178
rect -472 -186 -470 -178
rect -1167 -266 -1165 -258
rect -756 -262 -754 -254
rect -1240 -364 -1238 -356
rect -1174 -362 -1172 -354
rect -1146 -362 -1144 -354
rect -1077 -362 -1075 -354
rect -1049 -362 -1047 -354
rect -991 -362 -989 -354
rect -963 -362 -961 -354
rect -917 -362 -915 -354
rect -889 -362 -887 -354
rect -763 -362 -761 -354
rect -735 -362 -733 -354
rect -667 -362 -665 -354
rect -639 -362 -637 -354
rect -585 -362 -583 -354
rect -557 -362 -555 -354
rect -503 -362 -501 -354
rect -475 -362 -473 -354
rect -1170 -442 -1168 -434
rect -759 -438 -757 -430
rect -1232 -538 -1230 -530
rect -1166 -536 -1164 -528
rect -1138 -536 -1136 -528
rect -1069 -536 -1067 -528
rect -1041 -536 -1039 -528
rect -983 -536 -981 -528
rect -955 -536 -953 -528
rect -909 -536 -907 -528
rect -881 -536 -879 -528
rect -755 -536 -753 -528
rect -727 -536 -725 -528
rect -659 -536 -657 -528
rect -631 -536 -629 -528
rect -577 -536 -575 -528
rect -549 -536 -547 -528
rect -495 -536 -493 -528
rect -467 -536 -465 -528
rect -1162 -616 -1160 -608
rect -751 -612 -749 -604
<< polycontact >>
rect -1252 -22 -1248 -18
rect -1183 -18 -1179 -14
rect -1149 -18 -1145 -14
rect -1086 -18 -1082 -14
rect -1052 -18 -1048 -14
rect -1000 -18 -996 -14
rect -966 -18 -962 -14
rect -926 -18 -922 -14
rect -892 -18 -888 -14
rect -772 -18 -768 -14
rect -738 -18 -734 -14
rect -676 -18 -672 -14
rect -642 -18 -638 -14
rect -594 -18 -590 -14
rect -560 -18 -556 -14
rect -512 -18 -508 -14
rect -478 -18 -474 -14
rect -1182 -100 -1178 -96
rect -771 -96 -767 -92
rect -1244 -202 -1240 -198
rect -1175 -198 -1171 -194
rect -1141 -198 -1137 -194
rect -1078 -198 -1074 -194
rect -1044 -198 -1040 -194
rect -992 -198 -988 -194
rect -958 -198 -954 -194
rect -918 -198 -914 -194
rect -884 -198 -880 -194
rect -764 -198 -760 -194
rect -730 -198 -726 -194
rect -668 -198 -664 -194
rect -634 -198 -630 -194
rect -586 -198 -582 -194
rect -552 -198 -548 -194
rect -504 -198 -500 -194
rect -470 -198 -466 -194
rect -1174 -280 -1170 -276
rect -763 -276 -759 -272
rect -1247 -378 -1243 -374
rect -1178 -374 -1174 -370
rect -1144 -374 -1140 -370
rect -1081 -374 -1077 -370
rect -1047 -374 -1043 -370
rect -995 -374 -991 -370
rect -961 -374 -957 -370
rect -921 -374 -917 -370
rect -887 -374 -883 -370
rect -767 -374 -763 -370
rect -733 -374 -729 -370
rect -671 -374 -667 -370
rect -637 -374 -633 -370
rect -589 -374 -585 -370
rect -555 -374 -551 -370
rect -507 -374 -503 -370
rect -473 -374 -469 -370
rect -1177 -456 -1173 -452
rect -766 -452 -762 -448
rect -1239 -552 -1235 -548
rect -1170 -548 -1166 -544
rect -1136 -548 -1132 -544
rect -1073 -548 -1069 -544
rect -1039 -548 -1035 -544
rect -987 -548 -983 -544
rect -953 -548 -949 -544
rect -913 -548 -909 -544
rect -879 -548 -875 -544
rect -759 -548 -755 -544
rect -725 -548 -721 -544
rect -663 -548 -659 -544
rect -629 -548 -625 -544
rect -581 -548 -577 -544
rect -547 -548 -543 -544
rect -499 -548 -495 -544
rect -465 -548 -461 -544
rect -1169 -630 -1165 -626
rect -758 -626 -754 -622
<< ndcontact >>
rect -1252 -33 -1248 -28
rect -1240 -33 -1236 -28
rect -1186 -32 -1182 -27
rect -1174 -32 -1170 -27
rect -1158 -32 -1154 -27
rect -1146 -32 -1142 -27
rect -1089 -32 -1085 -27
rect -1077 -32 -1073 -27
rect -1061 -32 -1057 -27
rect -1049 -32 -1045 -27
rect -1003 -32 -999 -27
rect -991 -32 -987 -27
rect -975 -32 -971 -27
rect -963 -32 -959 -27
rect -929 -32 -925 -27
rect -917 -32 -913 -27
rect -901 -32 -897 -27
rect -889 -32 -885 -27
rect -775 -32 -771 -27
rect -763 -32 -759 -27
rect -747 -32 -743 -27
rect -735 -32 -731 -27
rect -679 -32 -675 -27
rect -667 -32 -663 -27
rect -651 -32 -647 -27
rect -639 -32 -635 -27
rect -597 -32 -593 -27
rect -585 -32 -581 -27
rect -569 -32 -565 -27
rect -557 -32 -553 -27
rect -515 -32 -511 -27
rect -503 -32 -499 -27
rect -487 -32 -483 -27
rect -475 -32 -471 -27
rect -1182 -111 -1178 -106
rect -1170 -111 -1166 -106
rect -771 -107 -767 -102
rect -759 -107 -755 -102
rect -1244 -213 -1240 -208
rect -1232 -213 -1228 -208
rect -1178 -212 -1174 -207
rect -1166 -212 -1162 -207
rect -1150 -212 -1146 -207
rect -1138 -212 -1134 -207
rect -1081 -212 -1077 -207
rect -1069 -212 -1065 -207
rect -1053 -212 -1049 -207
rect -1041 -212 -1037 -207
rect -995 -212 -991 -207
rect -983 -212 -979 -207
rect -967 -212 -963 -207
rect -955 -212 -951 -207
rect -921 -212 -917 -207
rect -909 -212 -905 -207
rect -893 -212 -889 -207
rect -881 -212 -877 -207
rect -767 -212 -763 -207
rect -755 -212 -751 -207
rect -739 -212 -735 -207
rect -727 -212 -723 -207
rect -671 -212 -667 -207
rect -659 -212 -655 -207
rect -643 -212 -639 -207
rect -631 -212 -627 -207
rect -589 -212 -585 -207
rect -577 -212 -573 -207
rect -561 -212 -557 -207
rect -549 -212 -545 -207
rect -507 -212 -503 -207
rect -495 -212 -491 -207
rect -479 -212 -475 -207
rect -467 -212 -463 -207
rect -1174 -291 -1170 -286
rect -1162 -291 -1158 -286
rect -763 -287 -759 -282
rect -751 -287 -747 -282
rect -1247 -389 -1243 -384
rect -1235 -389 -1231 -384
rect -1181 -388 -1177 -383
rect -1169 -388 -1165 -383
rect -1153 -388 -1149 -383
rect -1141 -388 -1137 -383
rect -1084 -388 -1080 -383
rect -1072 -388 -1068 -383
rect -1056 -388 -1052 -383
rect -1044 -388 -1040 -383
rect -998 -388 -994 -383
rect -986 -388 -982 -383
rect -970 -388 -966 -383
rect -958 -388 -954 -383
rect -924 -388 -920 -383
rect -912 -388 -908 -383
rect -896 -388 -892 -383
rect -884 -388 -880 -383
rect -770 -388 -766 -383
rect -758 -388 -754 -383
rect -742 -388 -738 -383
rect -730 -388 -726 -383
rect -674 -388 -670 -383
rect -662 -388 -658 -383
rect -646 -388 -642 -383
rect -634 -388 -630 -383
rect -592 -388 -588 -383
rect -580 -388 -576 -383
rect -564 -388 -560 -383
rect -552 -388 -548 -383
rect -510 -388 -506 -383
rect -498 -388 -494 -383
rect -482 -388 -478 -383
rect -470 -388 -466 -383
rect -1177 -467 -1173 -462
rect -1165 -467 -1161 -462
rect -766 -463 -762 -458
rect -754 -463 -750 -458
rect -1239 -563 -1235 -558
rect -1227 -563 -1223 -558
rect -1173 -562 -1169 -557
rect -1161 -562 -1157 -557
rect -1145 -562 -1141 -557
rect -1133 -562 -1129 -557
rect -1076 -562 -1072 -557
rect -1064 -562 -1060 -557
rect -1048 -562 -1044 -557
rect -1036 -562 -1032 -557
rect -990 -562 -986 -557
rect -978 -562 -974 -557
rect -962 -562 -958 -557
rect -950 -562 -946 -557
rect -916 -562 -912 -557
rect -904 -562 -900 -557
rect -888 -562 -884 -557
rect -876 -562 -872 -557
rect -762 -562 -758 -557
rect -750 -562 -746 -557
rect -734 -562 -730 -557
rect -722 -562 -718 -557
rect -666 -562 -662 -557
rect -654 -562 -650 -557
rect -638 -562 -634 -557
rect -626 -562 -622 -557
rect -584 -562 -580 -557
rect -572 -562 -568 -557
rect -556 -562 -552 -557
rect -544 -562 -540 -557
rect -502 -562 -498 -557
rect -490 -562 -486 -557
rect -474 -562 -470 -557
rect -462 -562 -458 -557
rect -1169 -641 -1165 -636
rect -1157 -641 -1153 -636
rect -758 -637 -754 -632
rect -746 -637 -742 -632
<< pdcontact >>
rect -1252 -8 -1248 0
rect -1240 -8 -1236 0
rect -1185 -6 -1181 2
rect -1175 -6 -1171 2
rect -1157 -6 -1153 2
rect -1147 -6 -1143 2
rect -1088 -6 -1084 2
rect -1078 -6 -1074 2
rect -1060 -6 -1056 2
rect -1050 -6 -1046 2
rect -1002 -6 -998 2
rect -992 -6 -988 2
rect -974 -6 -970 2
rect -964 -6 -960 2
rect -928 -6 -924 2
rect -918 -6 -914 2
rect -900 -6 -896 2
rect -890 -6 -886 2
rect -774 -6 -770 2
rect -764 -6 -760 2
rect -746 -6 -742 2
rect -736 -6 -732 2
rect -678 -6 -674 2
rect -668 -6 -664 2
rect -650 -6 -646 2
rect -640 -6 -636 2
rect -596 -6 -592 2
rect -586 -6 -582 2
rect -568 -6 -564 2
rect -558 -6 -554 2
rect -514 -6 -510 2
rect -504 -6 -500 2
rect -486 -6 -482 2
rect -476 -6 -472 2
rect -1182 -86 -1178 -78
rect -1170 -86 -1166 -78
rect -771 -82 -767 -74
rect -759 -82 -755 -74
rect -1244 -188 -1240 -180
rect -1232 -188 -1228 -180
rect -1177 -186 -1173 -178
rect -1167 -186 -1163 -178
rect -1149 -186 -1145 -178
rect -1139 -186 -1135 -178
rect -1080 -186 -1076 -178
rect -1070 -186 -1066 -178
rect -1052 -186 -1048 -178
rect -1042 -186 -1038 -178
rect -994 -186 -990 -178
rect -984 -186 -980 -178
rect -966 -186 -962 -178
rect -956 -186 -952 -178
rect -920 -186 -916 -178
rect -910 -186 -906 -178
rect -892 -186 -888 -178
rect -882 -186 -878 -178
rect -766 -186 -762 -178
rect -756 -186 -752 -178
rect -738 -186 -734 -178
rect -728 -186 -724 -178
rect -670 -186 -666 -178
rect -660 -186 -656 -178
rect -642 -186 -638 -178
rect -632 -186 -628 -178
rect -588 -186 -584 -178
rect -578 -186 -574 -178
rect -560 -186 -556 -178
rect -550 -186 -546 -178
rect -506 -186 -502 -178
rect -496 -186 -492 -178
rect -478 -186 -474 -178
rect -468 -186 -464 -178
rect -1174 -266 -1170 -258
rect -1162 -266 -1158 -258
rect -763 -262 -759 -254
rect -751 -262 -747 -254
rect -1247 -364 -1243 -356
rect -1235 -364 -1231 -356
rect -1180 -362 -1176 -354
rect -1170 -362 -1166 -354
rect -1152 -362 -1148 -354
rect -1142 -362 -1138 -354
rect -1083 -362 -1079 -354
rect -1073 -362 -1069 -354
rect -1055 -362 -1051 -354
rect -1045 -362 -1041 -354
rect -997 -362 -993 -354
rect -987 -362 -983 -354
rect -969 -362 -965 -354
rect -959 -362 -955 -354
rect -923 -362 -919 -354
rect -913 -362 -909 -354
rect -895 -362 -891 -354
rect -885 -362 -881 -354
rect -769 -362 -765 -354
rect -759 -362 -755 -354
rect -741 -362 -737 -354
rect -731 -362 -727 -354
rect -673 -362 -669 -354
rect -663 -362 -659 -354
rect -645 -362 -641 -354
rect -635 -362 -631 -354
rect -591 -362 -587 -354
rect -581 -362 -577 -354
rect -563 -362 -559 -354
rect -553 -362 -549 -354
rect -509 -362 -505 -354
rect -499 -362 -495 -354
rect -481 -362 -477 -354
rect -471 -362 -467 -354
rect -1177 -442 -1173 -434
rect -1165 -442 -1161 -434
rect -766 -438 -762 -430
rect -754 -438 -750 -430
rect -1239 -538 -1235 -530
rect -1227 -538 -1223 -530
rect -1172 -536 -1168 -528
rect -1162 -536 -1158 -528
rect -1144 -536 -1140 -528
rect -1134 -536 -1130 -528
rect -1075 -536 -1071 -528
rect -1065 -536 -1061 -528
rect -1047 -536 -1043 -528
rect -1037 -536 -1033 -528
rect -989 -536 -985 -528
rect -979 -536 -975 -528
rect -961 -536 -957 -528
rect -951 -536 -947 -528
rect -915 -536 -911 -528
rect -905 -536 -901 -528
rect -887 -536 -883 -528
rect -877 -536 -873 -528
rect -761 -536 -757 -528
rect -751 -536 -747 -528
rect -733 -536 -729 -528
rect -723 -536 -719 -528
rect -665 -536 -661 -528
rect -655 -536 -651 -528
rect -637 -536 -633 -528
rect -627 -536 -623 -528
rect -583 -536 -579 -528
rect -573 -536 -569 -528
rect -555 -536 -551 -528
rect -545 -536 -541 -528
rect -501 -536 -497 -528
rect -491 -536 -487 -528
rect -473 -536 -469 -528
rect -463 -536 -459 -528
rect -1169 -616 -1165 -608
rect -1157 -616 -1153 -608
rect -758 -612 -754 -604
rect -746 -612 -742 -604
<< m2contact >>
rect -1300 4 -1296 8
rect -1221 11 -1217 15
rect -833 4 -829 8
rect -869 -1 -864 4
rect -1270 -22 -1265 -18
rect -1125 -10 -1121 -6
rect -1104 -18 -1100 -14
rect -1028 -10 -1024 -6
rect -950 -10 -946 -6
rect -878 -18 -874 -14
rect -1118 -25 -1114 -21
rect -455 -1 -450 4
rect -714 -10 -710 -6
rect -694 -18 -690 -14
rect -618 -10 -614 -6
rect -536 -10 -532 -6
rect -464 -18 -460 -14
rect -1201 -40 -1197 -36
rect -706 -25 -702 -21
rect -790 -40 -786 -36
rect -1351 -124 -1347 -120
rect -1287 -59 -1282 -54
rect -1104 -55 -1100 -51
rect -1213 -65 -1209 -61
rect -1200 -73 -1196 -69
rect -694 -55 -690 -51
rect -802 -59 -798 -55
rect -789 -69 -785 -65
rect -1292 -176 -1288 -172
rect -1213 -169 -1209 -165
rect -825 -176 -821 -172
rect -861 -181 -856 -176
rect -1262 -202 -1257 -198
rect -1117 -190 -1113 -186
rect -1096 -198 -1092 -194
rect -1020 -190 -1016 -186
rect -942 -190 -938 -186
rect -870 -198 -866 -194
rect -1110 -205 -1106 -201
rect -447 -181 -442 -176
rect -706 -190 -702 -186
rect -686 -198 -682 -194
rect -610 -190 -606 -186
rect -528 -190 -524 -186
rect -456 -198 -452 -194
rect -1193 -220 -1189 -216
rect -1351 -228 -1347 -224
rect -698 -205 -694 -201
rect -423 -211 -419 -207
rect -782 -220 -778 -216
rect -1279 -239 -1274 -234
rect -1096 -235 -1092 -231
rect -1205 -245 -1201 -241
rect -1192 -253 -1188 -249
rect -686 -235 -682 -231
rect -794 -239 -790 -235
rect -781 -249 -777 -245
rect -1295 -352 -1291 -348
rect -1216 -345 -1212 -341
rect -828 -352 -824 -348
rect -864 -357 -859 -352
rect -1265 -378 -1260 -374
rect -1120 -366 -1116 -362
rect -1099 -374 -1095 -370
rect -1023 -366 -1019 -362
rect -945 -366 -941 -362
rect -873 -374 -869 -370
rect -1113 -381 -1109 -377
rect -450 -357 -445 -352
rect -709 -366 -705 -362
rect -689 -374 -685 -370
rect -613 -366 -609 -362
rect -531 -366 -527 -362
rect -459 -374 -455 -370
rect -1196 -396 -1192 -392
rect -1351 -404 -1347 -400
rect -701 -381 -697 -377
rect -425 -387 -421 -383
rect -785 -396 -781 -392
rect -1282 -415 -1277 -410
rect -1099 -411 -1095 -407
rect -1208 -421 -1204 -417
rect -1195 -429 -1191 -425
rect -689 -411 -685 -407
rect -797 -415 -793 -411
rect -784 -425 -780 -421
rect -1287 -526 -1283 -522
rect -1208 -519 -1204 -515
rect -820 -526 -816 -522
rect -856 -531 -851 -526
rect -1257 -552 -1252 -548
rect -1112 -540 -1108 -536
rect -1091 -548 -1087 -544
rect -1015 -540 -1011 -536
rect -937 -540 -933 -536
rect -865 -548 -861 -544
rect -1105 -555 -1101 -551
rect -442 -531 -437 -526
rect -701 -540 -697 -536
rect -681 -548 -677 -544
rect -605 -540 -601 -536
rect -523 -540 -519 -536
rect -451 -548 -447 -544
rect -1188 -570 -1184 -566
rect -1351 -578 -1347 -574
rect -693 -555 -689 -551
rect -417 -561 -413 -557
rect -777 -570 -773 -566
rect -1274 -589 -1269 -584
rect -1091 -585 -1087 -581
rect -1200 -595 -1196 -591
rect -1187 -603 -1183 -599
rect -681 -585 -677 -581
rect -789 -589 -785 -585
rect -776 -599 -772 -595
<< psubstratepcontact >>
rect -1252 -42 -1248 -38
rect -1146 -41 -1142 -37
rect -1049 -41 -1045 -37
rect -963 -41 -959 -37
rect -889 -41 -885 -37
rect -735 -41 -731 -37
rect -639 -41 -635 -37
rect -557 -41 -553 -37
rect -475 -41 -471 -37
rect -771 -116 -767 -112
rect -1182 -120 -1178 -116
rect -1244 -222 -1240 -218
rect -1138 -221 -1134 -217
rect -1041 -221 -1037 -217
rect -955 -221 -951 -217
rect -881 -221 -877 -217
rect -727 -221 -723 -217
rect -631 -221 -627 -217
rect -549 -221 -545 -217
rect -467 -221 -463 -217
rect -763 -296 -759 -292
rect -1174 -300 -1170 -296
rect -1247 -398 -1243 -394
rect -1141 -397 -1137 -393
rect -1044 -397 -1040 -393
rect -958 -397 -954 -393
rect -884 -397 -880 -393
rect -730 -397 -726 -393
rect -634 -397 -630 -393
rect -552 -397 -548 -393
rect -470 -397 -466 -393
rect -766 -472 -762 -468
rect -1177 -476 -1173 -472
rect -1239 -572 -1235 -568
rect -1133 -571 -1129 -567
rect -1036 -571 -1032 -567
rect -950 -571 -946 -567
rect -876 -571 -872 -567
rect -722 -571 -718 -567
rect -626 -571 -622 -567
rect -544 -571 -540 -567
rect -462 -571 -458 -567
rect -758 -646 -754 -642
rect -1169 -650 -1165 -646
<< nsubstratencontact >>
rect -1252 5 -1248 9
rect -1237 5 -1233 9
rect -1185 6 -1181 10
rect -1177 6 -1173 10
rect -1167 6 -1163 10
rect -1157 6 -1153 10
rect -1147 6 -1143 10
rect -1088 6 -1084 10
rect -1080 6 -1076 10
rect -1070 6 -1066 10
rect -1060 6 -1056 10
rect -1050 6 -1046 10
rect -1002 6 -998 10
rect -994 6 -990 10
rect -984 6 -980 10
rect -974 6 -970 10
rect -964 6 -960 10
rect -928 6 -924 10
rect -920 6 -916 10
rect -910 6 -906 10
rect -900 6 -896 10
rect -890 6 -886 10
rect -774 6 -770 10
rect -766 6 -762 10
rect -756 6 -752 10
rect -746 6 -742 10
rect -736 6 -732 10
rect -678 6 -674 10
rect -670 6 -666 10
rect -660 6 -656 10
rect -650 6 -646 10
rect -640 6 -636 10
rect -596 6 -592 10
rect -588 6 -584 10
rect -578 6 -574 10
rect -568 6 -564 10
rect -558 6 -554 10
rect -514 6 -510 10
rect -506 6 -502 10
rect -496 6 -492 10
rect -486 6 -482 10
rect -476 6 -472 10
rect -771 -69 -767 -65
rect -756 -69 -752 -65
rect -1182 -73 -1178 -69
rect -1167 -73 -1163 -69
rect -1244 -175 -1240 -171
rect -1229 -175 -1225 -171
rect -1177 -174 -1173 -170
rect -1169 -174 -1165 -170
rect -1159 -174 -1155 -170
rect -1149 -174 -1145 -170
rect -1139 -174 -1135 -170
rect -1080 -174 -1076 -170
rect -1072 -174 -1068 -170
rect -1062 -174 -1058 -170
rect -1052 -174 -1048 -170
rect -1042 -174 -1038 -170
rect -994 -174 -990 -170
rect -986 -174 -982 -170
rect -976 -174 -972 -170
rect -966 -174 -962 -170
rect -956 -174 -952 -170
rect -920 -174 -916 -170
rect -912 -174 -908 -170
rect -902 -174 -898 -170
rect -892 -174 -888 -170
rect -882 -174 -878 -170
rect -766 -174 -762 -170
rect -758 -174 -754 -170
rect -748 -174 -744 -170
rect -738 -174 -734 -170
rect -728 -174 -724 -170
rect -670 -174 -666 -170
rect -662 -174 -658 -170
rect -652 -174 -648 -170
rect -642 -174 -638 -170
rect -632 -174 -628 -170
rect -588 -174 -584 -170
rect -580 -174 -576 -170
rect -570 -174 -566 -170
rect -560 -174 -556 -170
rect -550 -174 -546 -170
rect -506 -174 -502 -170
rect -498 -174 -494 -170
rect -488 -174 -484 -170
rect -478 -174 -474 -170
rect -468 -174 -464 -170
rect -763 -249 -759 -245
rect -748 -249 -744 -245
rect -1174 -253 -1170 -249
rect -1159 -253 -1155 -249
rect -1247 -351 -1243 -347
rect -1232 -351 -1228 -347
rect -1180 -350 -1176 -346
rect -1172 -350 -1168 -346
rect -1162 -350 -1158 -346
rect -1152 -350 -1148 -346
rect -1142 -350 -1138 -346
rect -1083 -350 -1079 -346
rect -1075 -350 -1071 -346
rect -1065 -350 -1061 -346
rect -1055 -350 -1051 -346
rect -1045 -350 -1041 -346
rect -997 -350 -993 -346
rect -989 -350 -985 -346
rect -979 -350 -975 -346
rect -969 -350 -965 -346
rect -959 -350 -955 -346
rect -923 -350 -919 -346
rect -915 -350 -911 -346
rect -905 -350 -901 -346
rect -895 -350 -891 -346
rect -885 -350 -881 -346
rect -769 -350 -765 -346
rect -761 -350 -757 -346
rect -751 -350 -747 -346
rect -741 -350 -737 -346
rect -731 -350 -727 -346
rect -673 -350 -669 -346
rect -665 -350 -661 -346
rect -655 -350 -651 -346
rect -645 -350 -641 -346
rect -635 -350 -631 -346
rect -591 -350 -587 -346
rect -583 -350 -579 -346
rect -573 -350 -569 -346
rect -563 -350 -559 -346
rect -553 -350 -549 -346
rect -509 -350 -505 -346
rect -501 -350 -497 -346
rect -491 -350 -487 -346
rect -481 -350 -477 -346
rect -471 -350 -467 -346
rect -766 -425 -762 -421
rect -751 -425 -747 -421
rect -1177 -429 -1173 -425
rect -1162 -429 -1158 -425
rect -1239 -525 -1235 -521
rect -1224 -525 -1220 -521
rect -1172 -524 -1168 -520
rect -1164 -524 -1160 -520
rect -1154 -524 -1150 -520
rect -1144 -524 -1140 -520
rect -1134 -524 -1130 -520
rect -1075 -524 -1071 -520
rect -1067 -524 -1063 -520
rect -1057 -524 -1053 -520
rect -1047 -524 -1043 -520
rect -1037 -524 -1033 -520
rect -989 -524 -985 -520
rect -981 -524 -977 -520
rect -971 -524 -967 -520
rect -961 -524 -957 -520
rect -951 -524 -947 -520
rect -915 -524 -911 -520
rect -907 -524 -903 -520
rect -897 -524 -893 -520
rect -887 -524 -883 -520
rect -877 -524 -873 -520
rect -761 -524 -757 -520
rect -753 -524 -749 -520
rect -743 -524 -739 -520
rect -733 -524 -729 -520
rect -723 -524 -719 -520
rect -665 -524 -661 -520
rect -657 -524 -653 -520
rect -647 -524 -643 -520
rect -637 -524 -633 -520
rect -627 -524 -623 -520
rect -583 -524 -579 -520
rect -575 -524 -571 -520
rect -565 -524 -561 -520
rect -555 -524 -551 -520
rect -545 -524 -541 -520
rect -501 -524 -497 -520
rect -493 -524 -489 -520
rect -483 -524 -479 -520
rect -473 -524 -469 -520
rect -463 -524 -459 -520
rect -758 -599 -754 -595
rect -743 -599 -739 -595
rect -1169 -603 -1165 -599
rect -1154 -603 -1150 -599
<< labels >>
rlabel m2contact -1221 15 -1217 15 1 invout
rlabel metal1 -1236 -22 -1236 -17 1 invout
rlabel pdcontact -1185 1 -1185 1 1 M6source
rlabel pdcontact -1145 0 -1145 0 1 M7source
rlabel pdcontact -1088 1 -1088 1 1 M6source
rlabel pdcontact -1048 0 -1048 0 1 M7source
rlabel pdcontact -1002 1 -1002 1 1 M6source
rlabel pdcontact -962 0 -962 0 1 M7source
rlabel pdcontact -928 1 -928 1 1 M6source
rlabel pdcontact -888 0 -888 0 1 M7source
rlabel pdcontact -774 1 -774 1 1 M6source
rlabel pdcontact -734 0 -734 0 1 M7source
rlabel pdcontact -678 1 -678 1 1 M6source
rlabel pdcontact -638 0 -638 0 1 M7source
rlabel pdcontact -596 1 -596 1 1 M6source
rlabel pdcontact -556 0 -556 0 1 M7source
rlabel pdcontact -514 1 -514 1 1 M6source
rlabel pdcontact -474 0 -474 0 1 M7source
rlabel m2contact -1213 -165 -1209 -165 1 invout
rlabel metal1 -1228 -202 -1228 -197 1 invout
rlabel pdcontact -1177 -179 -1177 -179 1 M6source
rlabel pdcontact -1137 -180 -1137 -180 1 M7source
rlabel pdcontact -1080 -179 -1080 -179 1 M6source
rlabel pdcontact -1040 -180 -1040 -180 1 M7source
rlabel pdcontact -994 -179 -994 -179 1 M6source
rlabel pdcontact -954 -180 -954 -180 1 M7source
rlabel pdcontact -920 -179 -920 -179 1 M6source
rlabel pdcontact -880 -180 -880 -180 1 M7source
rlabel pdcontact -766 -179 -766 -179 1 M6source
rlabel pdcontact -726 -180 -726 -180 1 M7source
rlabel pdcontact -670 -179 -670 -179 1 M6source
rlabel pdcontact -630 -180 -630 -180 1 M7source
rlabel pdcontact -588 -179 -588 -179 1 M6source
rlabel pdcontact -548 -180 -548 -180 1 M7source
rlabel pdcontact -506 -179 -506 -179 1 M6source
rlabel pdcontact -466 -180 -466 -180 1 M7source
rlabel pdcontact -469 -356 -469 -356 1 M7source
rlabel pdcontact -509 -355 -509 -355 1 M6source
rlabel pdcontact -551 -356 -551 -356 1 M7source
rlabel pdcontact -591 -355 -591 -355 1 M6source
rlabel pdcontact -633 -356 -633 -356 1 M7source
rlabel pdcontact -673 -355 -673 -355 1 M6source
rlabel pdcontact -729 -356 -729 -356 1 M7source
rlabel pdcontact -769 -355 -769 -355 1 M6source
rlabel pdcontact -883 -356 -883 -356 1 M7source
rlabel pdcontact -923 -355 -923 -355 1 M6source
rlabel pdcontact -957 -356 -957 -356 1 M7source
rlabel pdcontact -997 -355 -997 -355 1 M6source
rlabel pdcontact -1043 -356 -1043 -356 1 M7source
rlabel pdcontact -1083 -355 -1083 -355 1 M6source
rlabel pdcontact -1140 -356 -1140 -356 1 M7source
rlabel pdcontact -1180 -355 -1180 -355 1 M6source
rlabel metal1 -1231 -378 -1231 -373 1 invout
rlabel m2contact -1216 -341 -1212 -341 1 invout
rlabel metal1 -1304 -589 -1304 -584 3 D
rlabel pdcontact -461 -530 -461 -530 1 M7source
rlabel pdcontact -501 -529 -501 -529 1 M6source
rlabel pdcontact -543 -530 -543 -530 1 M7source
rlabel pdcontact -583 -529 -583 -529 1 M6source
rlabel pdcontact -625 -530 -625 -530 1 M7source
rlabel pdcontact -665 -529 -665 -529 1 M6source
rlabel pdcontact -721 -530 -721 -530 1 M7source
rlabel pdcontact -761 -529 -761 -529 1 M6source
rlabel pdcontact -875 -530 -875 -530 1 M7source
rlabel pdcontact -915 -529 -915 -529 1 M6source
rlabel pdcontact -949 -530 -949 -530 1 M7source
rlabel pdcontact -989 -529 -989 -529 1 M6source
rlabel pdcontact -1035 -530 -1035 -530 1 M7source
rlabel pdcontact -1075 -529 -1075 -529 1 M6source
rlabel pdcontact -1132 -530 -1132 -530 1 M7source
rlabel pdcontact -1172 -529 -1172 -529 1 M6source
rlabel metal1 -1223 -552 -1223 -547 1 invout
rlabel m2contact -1208 -515 -1204 -515 1 invout
rlabel metal2 -1333 -670 -1330 -670 2 clock
rlabel metal1 -1362 -669 -1359 -669 2 vdd!
rlabel metal2 -1351 -668 -1347 -668 1 gnd!
<< end >>
