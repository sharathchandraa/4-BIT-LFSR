magic
tech scmos
timestamp 1398369974
<< nwell >>
rect -685 -12 -632 13
rect -549 -12 -496 13
rect -444 -12 -391 13
rect -347 -12 -294 13
rect -155 -10 -127 15
rect -87 -7 -34 18
rect 49 -7 102 18
rect 135 -7 188 18
rect 226 -7 279 18
rect -683 -106 -655 -81
rect -85 -101 -57 -76
<< polysilicon >>
rect -76 7 -74 9
rect -48 7 -46 9
rect 60 7 62 9
rect 88 7 90 9
rect 146 7 148 9
rect 174 7 176 9
rect 237 7 239 9
rect 265 7 267 9
rect -142 5 -140 7
rect -674 2 -672 4
rect -646 2 -644 4
rect -538 2 -536 4
rect -510 2 -508 4
rect -433 2 -431 4
rect -405 2 -403 4
rect -336 2 -334 4
rect -308 2 -306 4
rect -674 -27 -672 -6
rect -646 -27 -644 -6
rect -538 -27 -536 -6
rect -510 -27 -508 -6
rect -433 -27 -431 -6
rect -405 -27 -403 -6
rect -336 -27 -334 -6
rect -308 -27 -306 -6
rect -142 -14 -140 -3
rect -145 -16 -140 -14
rect -674 -33 -672 -31
rect -646 -33 -644 -31
rect -538 -33 -536 -31
rect -510 -33 -508 -31
rect -433 -33 -431 -31
rect -405 -33 -403 -31
rect -336 -33 -334 -31
rect -308 -33 -306 -31
rect -142 -24 -140 -16
rect -76 -22 -74 -1
rect -48 -22 -46 -1
rect 60 -22 62 -1
rect 88 -22 90 -1
rect 146 -22 148 -1
rect 174 -22 176 -1
rect 237 -22 239 -1
rect 265 -22 267 -1
rect -76 -28 -74 -26
rect -48 -28 -46 -26
rect 60 -28 62 -26
rect 88 -28 90 -26
rect 146 -28 148 -26
rect 174 -28 176 -26
rect 237 -28 239 -26
rect 265 -28 267 -26
rect -142 -30 -140 -28
rect -72 -86 -70 -84
rect -670 -91 -668 -89
rect -670 -110 -668 -99
rect -72 -105 -70 -94
rect -75 -107 -70 -105
rect -673 -112 -668 -110
rect -670 -120 -668 -112
rect -72 -115 -70 -107
rect -72 -121 -70 -119
rect -670 -126 -668 -124
<< ndiffusion >>
rect -677 -31 -674 -27
rect -672 -31 -669 -27
rect -649 -31 -646 -27
rect -644 -31 -641 -27
rect -541 -31 -538 -27
rect -536 -31 -533 -27
rect -513 -31 -510 -27
rect -508 -31 -505 -27
rect -436 -31 -433 -27
rect -431 -31 -428 -27
rect -408 -31 -405 -27
rect -403 -31 -400 -27
rect -339 -31 -336 -27
rect -334 -31 -331 -27
rect -311 -31 -308 -27
rect -306 -31 -303 -27
rect -145 -28 -142 -24
rect -140 -28 -137 -24
rect -79 -26 -76 -22
rect -74 -26 -71 -22
rect -51 -26 -48 -22
rect -46 -26 -43 -22
rect 57 -26 60 -22
rect 62 -26 65 -22
rect 85 -26 88 -22
rect 90 -26 93 -22
rect 143 -26 146 -22
rect 148 -26 151 -22
rect 171 -26 174 -22
rect 176 -26 179 -22
rect 234 -26 237 -22
rect 239 -26 242 -22
rect 262 -26 265 -22
rect 267 -26 270 -22
rect -75 -119 -72 -115
rect -70 -119 -67 -115
rect -673 -124 -670 -120
rect -668 -124 -665 -120
<< pdiffusion >>
rect -676 -6 -674 2
rect -672 -6 -670 2
rect -648 -6 -646 2
rect -644 -6 -642 2
rect -540 -6 -538 2
rect -536 -6 -534 2
rect -512 -6 -510 2
rect -508 -6 -506 2
rect -435 -6 -433 2
rect -431 -6 -429 2
rect -407 -6 -405 2
rect -403 -6 -401 2
rect -338 -6 -336 2
rect -334 -6 -332 2
rect -310 -6 -308 2
rect -306 -6 -304 2
rect -145 -3 -142 5
rect -140 -3 -137 5
rect -78 -1 -76 7
rect -74 -1 -72 7
rect -50 -1 -48 7
rect -46 -1 -44 7
rect 58 -1 60 7
rect 62 -1 64 7
rect 86 -1 88 7
rect 90 -1 92 7
rect 144 -1 146 7
rect 148 -1 150 7
rect 172 -1 174 7
rect 176 -1 178 7
rect 235 -1 237 7
rect 239 -1 241 7
rect 263 -1 265 7
rect 267 -1 269 7
rect -673 -99 -670 -91
rect -668 -99 -665 -91
rect -75 -94 -72 -86
rect -70 -94 -67 -86
<< metal1 >>
rect -236 25 253 28
rect -236 23 -232 25
rect -822 20 -232 23
rect -795 8 -791 20
rect -662 10 -658 20
rect -526 10 -522 20
rect -421 10 -417 20
rect -324 10 -320 20
rect -197 13 -193 25
rect -134 14 -130 25
rect -676 6 -672 10
rect -668 6 -662 10
rect -658 6 -652 10
rect -648 6 -642 10
rect -680 2 -676 6
rect -642 2 -638 6
rect -666 -6 -652 2
rect -540 6 -536 10
rect -532 6 -526 10
rect -522 6 -516 10
rect -512 6 -506 10
rect -544 2 -540 6
rect -506 2 -502 6
rect -530 -6 -516 2
rect -435 6 -431 10
rect -427 6 -421 10
rect -417 6 -411 10
rect -407 6 -401 10
rect -439 2 -435 6
rect -401 2 -397 6
rect -425 -6 -411 2
rect -338 6 -334 10
rect -330 6 -324 10
rect -320 6 -314 10
rect -310 6 -304 10
rect -145 10 -134 14
rect -342 2 -338 6
rect -304 2 -300 6
rect -149 5 -145 10
rect -328 -6 -314 2
rect -696 -18 -678 -14
rect -696 -36 -692 -18
rect -661 -21 -658 -6
rect -620 -14 -616 -10
rect -640 -18 -616 -14
rect -568 -18 -542 -14
rect -525 -21 -522 -6
rect -484 -14 -480 -10
rect -504 -18 -480 -14
rect -454 -18 -437 -14
rect -454 -21 -451 -18
rect -420 -21 -417 -6
rect -379 -14 -375 -10
rect -399 -18 -375 -14
rect -361 -18 -340 -14
rect -361 -21 -358 -18
rect -323 -21 -320 -6
rect -302 -18 -292 -14
rect -681 -24 -600 -21
rect -681 -27 -677 -24
rect -545 -24 -451 -21
rect -440 -24 -358 -21
rect -343 -24 -292 -21
rect -545 -27 -541 -24
rect -440 -27 -436 -24
rect -343 -27 -339 -24
rect -665 -32 -653 -27
rect -529 -32 -517 -27
rect -424 -32 -412 -27
rect -327 -32 -315 -27
rect -295 -28 -292 -24
rect -283 -27 -278 -1
rect -137 -13 -133 -3
rect -118 -13 -114 16
rect -64 15 -60 25
rect 72 15 76 25
rect 158 15 162 25
rect 249 15 253 25
rect -78 11 -74 15
rect -70 11 -64 15
rect -60 11 -54 15
rect -50 11 -44 15
rect -82 7 -78 11
rect -44 7 -40 11
rect -68 -1 -54 7
rect 58 11 62 15
rect 66 11 72 15
rect 76 11 82 15
rect 86 11 92 15
rect 54 7 58 11
rect 92 7 96 11
rect 68 -1 82 7
rect 144 11 148 15
rect 152 11 158 15
rect 162 11 168 15
rect 172 11 178 15
rect 140 7 144 11
rect 178 7 182 11
rect 154 -1 168 7
rect 235 11 239 15
rect 243 11 249 15
rect 253 11 259 15
rect 263 11 269 15
rect 231 7 235 11
rect 269 7 273 11
rect 245 -1 259 7
rect -162 -17 -149 -13
rect -137 -17 -114 -13
rect -98 -13 -80 -9
rect -137 -23 -133 -17
rect -283 -28 -218 -27
rect -295 -31 -218 -28
rect -641 -37 -637 -32
rect -641 -45 -637 -41
rect -505 -37 -501 -32
rect -505 -45 -501 -41
rect -400 -37 -396 -32
rect -400 -45 -396 -41
rect -303 -37 -299 -32
rect -149 -33 -145 -28
rect -98 -31 -94 -13
rect -63 -16 -60 -1
rect -22 -9 -18 -5
rect -42 -13 -18 -9
rect 30 -13 56 -9
rect 73 -16 76 -1
rect 114 -9 118 -5
rect 94 -13 118 -9
rect 125 -13 142 -9
rect 125 -16 128 -13
rect 159 -16 162 -1
rect 200 -9 204 -5
rect 180 -13 204 -9
rect 212 -13 233 -9
rect 212 -16 215 -13
rect 250 -16 253 -1
rect 271 -13 281 -9
rect -83 -19 -2 -16
rect -83 -22 -79 -19
rect 53 -19 128 -16
rect 139 -19 215 -16
rect 230 -19 281 -16
rect 53 -22 57 -19
rect 139 -22 143 -19
rect 230 -22 234 -19
rect -67 -27 -55 -22
rect 69 -27 81 -22
rect 155 -27 167 -22
rect 246 -27 258 -22
rect 278 -23 281 -19
rect 290 -23 295 4
rect 278 -26 303 -23
rect -43 -32 -39 -27
rect -149 -40 -145 -37
rect -43 -40 -39 -36
rect 93 -32 97 -27
rect 93 -40 97 -36
rect 179 -32 183 -27
rect 179 -40 183 -36
rect 270 -32 274 -27
rect 270 -40 274 -36
rect -303 -45 -299 -41
rect -230 -43 274 -40
rect -230 -45 -225 -43
rect -809 -48 -225 -45
rect -816 -59 -782 -54
rect -729 -136 -725 -48
rect -214 -54 -184 -49
rect -708 -109 -704 -69
rect -691 -86 -677 -82
rect -673 -86 -662 -82
rect -677 -91 -673 -86
rect -665 -109 -661 -99
rect -572 -109 -568 -65
rect -708 -113 -677 -109
rect -665 -113 -568 -109
rect -665 -119 -661 -113
rect -677 -129 -673 -124
rect -677 -136 -673 -133
rect -131 -131 -127 -43
rect -110 -104 -106 -64
rect -93 -81 -79 -77
rect -75 -81 -64 -77
rect -79 -86 -75 -81
rect -67 -104 -63 -94
rect 26 -104 30 -60
rect -110 -108 -79 -104
rect -67 -108 30 -104
rect -67 -114 -63 -108
rect -79 -124 -75 -119
rect -79 -131 -75 -128
rect -131 -134 -75 -131
rect -729 -139 -673 -136
<< metal2 >>
rect -484 86 -480 87
rect -484 81 -162 86
rect -484 36 -480 81
rect -831 33 -480 36
rect -795 -82 -791 4
rect -620 -6 -616 33
rect -484 -6 -480 33
rect -379 31 -278 35
rect -379 -6 -375 31
rect -283 4 -278 31
rect -288 -18 -246 -14
rect -708 -40 -696 -36
rect -708 -54 -704 -40
rect -777 -59 -704 -54
rect -708 -65 -704 -59
rect -600 -79 -596 -25
rect -572 -61 -568 -18
rect -252 -79 -246 -18
rect -218 -49 -214 -31
rect -600 -82 -246 -79
rect -197 -77 -193 9
rect -167 -13 -162 81
rect -118 38 118 41
rect -118 20 -114 38
rect -22 -1 -18 38
rect 114 -1 118 38
rect 200 36 295 40
rect 200 -1 204 36
rect 290 9 295 36
rect 285 -13 314 -9
rect -110 -35 -98 -31
rect -110 -49 -106 -35
rect -179 -54 -106 -49
rect -110 -60 -106 -54
rect -2 -74 2 -20
rect 26 -56 30 -13
rect 308 -74 314 -13
rect -2 -77 314 -74
rect -197 -81 -97 -77
rect -1 -78 314 -77
rect -795 -86 -695 -82
rect -599 -83 -246 -82
<< ntransistor >>
rect -674 -31 -672 -27
rect -646 -31 -644 -27
rect -538 -31 -536 -27
rect -510 -31 -508 -27
rect -433 -31 -431 -27
rect -405 -31 -403 -27
rect -336 -31 -334 -27
rect -308 -31 -306 -27
rect -142 -28 -140 -24
rect -76 -26 -74 -22
rect -48 -26 -46 -22
rect 60 -26 62 -22
rect 88 -26 90 -22
rect 146 -26 148 -22
rect 174 -26 176 -22
rect 237 -26 239 -22
rect 265 -26 267 -22
rect -72 -119 -70 -115
rect -670 -124 -668 -120
<< ptransistor >>
rect -674 -6 -672 2
rect -646 -6 -644 2
rect -538 -6 -536 2
rect -510 -6 -508 2
rect -433 -6 -431 2
rect -405 -6 -403 2
rect -336 -6 -334 2
rect -308 -6 -306 2
rect -142 -3 -140 5
rect -76 -1 -74 7
rect -48 -1 -46 7
rect 60 -1 62 7
rect 88 -1 90 7
rect 146 -1 148 7
rect 174 -1 176 7
rect 237 -1 239 7
rect 265 -1 267 7
rect -670 -99 -668 -91
rect -72 -94 -70 -86
<< polycontact >>
rect -678 -18 -674 -14
rect -644 -18 -640 -14
rect -542 -18 -538 -14
rect -508 -18 -504 -14
rect -437 -18 -433 -14
rect -403 -18 -399 -14
rect -340 -18 -336 -14
rect -306 -18 -302 -14
rect -149 -17 -145 -13
rect -80 -13 -76 -9
rect -46 -13 -42 -9
rect 56 -13 60 -9
rect 90 -13 94 -9
rect 142 -13 146 -9
rect 176 -13 180 -9
rect 233 -13 237 -9
rect 267 -13 271 -9
rect -677 -113 -673 -109
rect -79 -108 -75 -104
<< ndcontact >>
rect -681 -32 -677 -27
rect -669 -32 -665 -27
rect -653 -32 -649 -27
rect -641 -32 -637 -27
rect -545 -32 -541 -27
rect -533 -32 -529 -27
rect -517 -32 -513 -27
rect -505 -32 -501 -27
rect -440 -32 -436 -27
rect -428 -32 -424 -27
rect -412 -32 -408 -27
rect -400 -32 -396 -27
rect -343 -32 -339 -27
rect -331 -32 -327 -27
rect -315 -32 -311 -27
rect -303 -32 -299 -27
rect -149 -28 -145 -23
rect -137 -28 -133 -23
rect -83 -27 -79 -22
rect -71 -27 -67 -22
rect -55 -27 -51 -22
rect -43 -27 -39 -22
rect 53 -27 57 -22
rect 65 -27 69 -22
rect 81 -27 85 -22
rect 93 -27 97 -22
rect 139 -27 143 -22
rect 151 -27 155 -22
rect 167 -27 171 -22
rect 179 -27 183 -22
rect 230 -27 234 -22
rect 242 -27 246 -22
rect 258 -27 262 -22
rect 270 -27 274 -22
rect -677 -124 -673 -119
rect -79 -119 -75 -114
rect -67 -119 -63 -114
rect -665 -124 -661 -119
<< pdcontact >>
rect -680 -6 -676 2
rect -670 -6 -666 2
rect -652 -6 -648 2
rect -642 -6 -638 2
rect -544 -6 -540 2
rect -534 -6 -530 2
rect -516 -6 -512 2
rect -506 -6 -502 2
rect -439 -6 -435 2
rect -429 -6 -425 2
rect -411 -6 -407 2
rect -401 -6 -397 2
rect -342 -6 -338 2
rect -332 -6 -328 2
rect -314 -6 -310 2
rect -304 -6 -300 2
rect -149 -3 -145 5
rect -137 -3 -133 5
rect -82 -1 -78 7
rect -72 -1 -68 7
rect -54 -1 -50 7
rect -44 -1 -40 7
rect 54 -1 58 7
rect 64 -1 68 7
rect 82 -1 86 7
rect 92 -1 96 7
rect 140 -1 144 7
rect 150 -1 154 7
rect 168 -1 172 7
rect 178 -1 182 7
rect 231 -1 235 7
rect 241 -1 245 7
rect 259 -1 263 7
rect 269 -1 273 7
rect -677 -99 -673 -91
rect -665 -99 -661 -91
rect -79 -94 -75 -86
rect -67 -94 -63 -86
<< m2contact >>
rect -795 4 -791 8
rect -197 9 -193 13
rect -118 16 -114 20
rect -283 -1 -278 4
rect -620 -10 -616 -6
rect -572 -18 -568 -14
rect -484 -10 -480 -6
rect -379 -10 -375 -6
rect -292 -18 -288 -14
rect -600 -25 -596 -21
rect 290 4 295 9
rect -167 -17 -162 -13
rect -218 -31 -214 -27
rect -696 -40 -692 -36
rect -22 -5 -18 -1
rect 26 -13 30 -9
rect 114 -5 118 -1
rect 200 -5 204 -1
rect 281 -13 285 -9
rect -2 -20 2 -16
rect -98 -35 -94 -31
rect -782 -59 -777 -54
rect -218 -54 -214 -49
rect -184 -54 -179 -49
rect -572 -65 -568 -61
rect -708 -69 -704 -65
rect -695 -86 -691 -82
rect 26 -60 30 -56
rect -110 -64 -106 -60
rect -97 -81 -93 -77
<< psubstratepcontact >>
rect -149 -37 -145 -33
rect -43 -36 -39 -32
rect 93 -36 97 -32
rect 179 -36 183 -32
rect 270 -36 274 -32
rect -641 -41 -637 -37
rect -505 -41 -501 -37
rect -400 -41 -396 -37
rect -303 -41 -299 -37
rect -79 -128 -75 -124
rect -677 -133 -673 -129
<< nsubstratencontact >>
rect -149 10 -145 14
rect -134 10 -130 14
rect -82 11 -78 15
rect -74 11 -70 15
rect -64 11 -60 15
rect -54 11 -50 15
rect -44 11 -40 15
rect 54 11 58 15
rect 62 11 66 15
rect 72 11 76 15
rect 82 11 86 15
rect 92 11 96 15
rect 140 11 144 15
rect 148 11 152 15
rect 158 11 162 15
rect 168 11 172 15
rect 178 11 182 15
rect 231 11 235 15
rect 239 11 243 15
rect 249 11 253 15
rect 259 11 263 15
rect 269 11 273 15
rect -680 6 -676 10
rect -672 6 -668 10
rect -662 6 -658 10
rect -652 6 -648 10
rect -642 6 -638 10
rect -544 6 -540 10
rect -536 6 -532 10
rect -526 6 -522 10
rect -516 6 -512 10
rect -506 6 -502 10
rect -439 6 -435 10
rect -431 6 -427 10
rect -421 6 -417 10
rect -411 6 -407 10
rect -401 6 -397 10
rect -342 6 -338 10
rect -334 6 -330 10
rect -324 6 -320 10
rect -314 6 -310 10
rect -304 6 -300 10
rect -79 -81 -75 -77
rect -64 -81 -60 -77
rect -677 -86 -673 -82
rect -662 -86 -658 -82
<< labels >>
rlabel pdcontact -439 1 -439 1 1 M6source
rlabel pdcontact -399 0 -399 0 1 M7source
rlabel pdcontact -680 1 -680 1 1 M6source
rlabel pdcontact -640 0 -640 0 1 M7source
rlabel pdcontact -544 1 -544 1 1 M6source
rlabel pdcontact -504 0 -504 0 1 M7source
rlabel metal1 -822 20 -822 23 3 vdd!
rlabel metal1 -809 -48 -809 -45 1 gnd!
rlabel metal1 -816 -59 -816 -54 1 D
rlabel metal2 -831 33 -831 36 3 clock
rlabel pdcontact -342 1 -342 1 1 M6source
rlabel pdcontact -302 0 -302 0 1 M7source
rlabel m2contact -118 20 -114 20 1 invout
rlabel metal1 -133 -17 -133 -12 1 invout
rlabel pdcontact -82 6 -82 6 1 M6source
rlabel pdcontact -42 5 -42 5 1 M7source
rlabel pdcontact 54 6 54 6 1 M6source
rlabel pdcontact 94 5 94 5 1 M7source
rlabel pdcontact 140 6 140 6 1 M6source
rlabel pdcontact 180 5 180 5 1 M7source
rlabel pdcontact 231 6 231 6 1 M6source
rlabel pdcontact 271 5 271 5 1 M7source
rlabel metal1 303 -26 303 -23 7 Q
<< end >>
