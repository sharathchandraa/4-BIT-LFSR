magic
tech scmos
timestamp 1398571937
<< nwell >>
rect -1258 -15 -1230 10
rect -1190 -12 -1137 13
rect -1093 -12 -1040 13
rect -1007 -12 -954 13
rect -933 -12 -880 13
rect -779 -12 -726 13
rect -683 -12 -630 13
rect -601 -12 -548 13
rect -519 -12 -466 13
rect -1188 -93 -1160 -68
rect -777 -89 -749 -64
<< polysilicon >>
rect -1179 2 -1177 4
rect -1151 2 -1149 4
rect -1082 2 -1080 4
rect -1054 2 -1052 4
rect -996 2 -994 4
rect -968 2 -966 4
rect -922 2 -920 4
rect -894 2 -892 4
rect -768 2 -766 4
rect -740 2 -738 4
rect -672 2 -670 4
rect -644 2 -642 4
rect -590 2 -588 4
rect -562 2 -560 4
rect -508 2 -506 4
rect -480 2 -478 4
rect -1245 0 -1243 2
rect -1245 -19 -1243 -8
rect -1248 -21 -1243 -19
rect -1245 -29 -1243 -21
rect -1179 -27 -1177 -6
rect -1151 -27 -1149 -6
rect -1082 -27 -1080 -6
rect -1054 -27 -1052 -6
rect -996 -27 -994 -6
rect -968 -27 -966 -6
rect -922 -27 -920 -6
rect -894 -27 -892 -6
rect -768 -27 -766 -6
rect -740 -27 -738 -6
rect -672 -27 -670 -6
rect -644 -27 -642 -6
rect -590 -27 -588 -6
rect -562 -27 -560 -6
rect -508 -27 -506 -6
rect -480 -27 -478 -6
rect -1179 -33 -1177 -31
rect -1151 -33 -1149 -31
rect -1082 -33 -1080 -31
rect -1054 -33 -1052 -31
rect -996 -33 -994 -31
rect -968 -33 -966 -31
rect -922 -33 -920 -31
rect -894 -33 -892 -31
rect -768 -33 -766 -31
rect -740 -33 -738 -31
rect -672 -33 -670 -31
rect -644 -33 -642 -31
rect -590 -33 -588 -31
rect -562 -33 -560 -31
rect -508 -33 -506 -31
rect -480 -33 -478 -31
rect -1245 -35 -1243 -33
rect -764 -74 -762 -72
rect -1175 -78 -1173 -76
rect -1175 -97 -1173 -86
rect -764 -93 -762 -82
rect -767 -95 -762 -93
rect -1178 -99 -1173 -97
rect -1175 -107 -1173 -99
rect -764 -103 -762 -95
rect -764 -109 -762 -107
rect -1175 -113 -1173 -111
<< ndiffusion >>
rect -1248 -33 -1245 -29
rect -1243 -33 -1240 -29
rect -1182 -31 -1179 -27
rect -1177 -31 -1174 -27
rect -1154 -31 -1151 -27
rect -1149 -31 -1146 -27
rect -1085 -31 -1082 -27
rect -1080 -31 -1077 -27
rect -1057 -31 -1054 -27
rect -1052 -31 -1049 -27
rect -999 -31 -996 -27
rect -994 -31 -991 -27
rect -971 -31 -968 -27
rect -966 -31 -963 -27
rect -925 -31 -922 -27
rect -920 -31 -917 -27
rect -897 -31 -894 -27
rect -892 -31 -889 -27
rect -771 -31 -768 -27
rect -766 -31 -763 -27
rect -743 -31 -740 -27
rect -738 -31 -735 -27
rect -675 -31 -672 -27
rect -670 -31 -667 -27
rect -647 -31 -644 -27
rect -642 -31 -639 -27
rect -593 -31 -590 -27
rect -588 -31 -585 -27
rect -565 -31 -562 -27
rect -560 -31 -557 -27
rect -511 -31 -508 -27
rect -506 -31 -503 -27
rect -483 -31 -480 -27
rect -478 -31 -475 -27
rect -1178 -111 -1175 -107
rect -1173 -111 -1170 -107
rect -767 -107 -764 -103
rect -762 -107 -759 -103
<< pdiffusion >>
rect -1248 -8 -1245 0
rect -1243 -8 -1240 0
rect -1181 -6 -1179 2
rect -1177 -6 -1175 2
rect -1153 -6 -1151 2
rect -1149 -6 -1147 2
rect -1084 -6 -1082 2
rect -1080 -6 -1078 2
rect -1056 -6 -1054 2
rect -1052 -6 -1050 2
rect -998 -6 -996 2
rect -994 -6 -992 2
rect -970 -6 -968 2
rect -966 -6 -964 2
rect -924 -6 -922 2
rect -920 -6 -918 2
rect -896 -6 -894 2
rect -892 -6 -890 2
rect -770 -6 -768 2
rect -766 -6 -764 2
rect -742 -6 -740 2
rect -738 -6 -736 2
rect -674 -6 -672 2
rect -670 -6 -668 2
rect -646 -6 -644 2
rect -642 -6 -640 2
rect -592 -6 -590 2
rect -588 -6 -586 2
rect -564 -6 -562 2
rect -560 -6 -558 2
rect -510 -6 -508 2
rect -506 -6 -504 2
rect -482 -6 -480 2
rect -478 -6 -476 2
rect -1178 -86 -1175 -78
rect -1173 -86 -1170 -78
rect -767 -82 -764 -74
rect -762 -82 -759 -74
<< metal1 >>
rect -1311 20 -492 23
rect -1300 8 -1296 20
rect -1237 9 -1233 20
rect -1248 5 -1237 9
rect -1252 0 -1248 5
rect -1240 -18 -1236 -8
rect -1221 -18 -1217 11
rect -1167 10 -1163 20
rect -1070 10 -1066 20
rect -984 10 -980 20
rect -910 10 -906 20
rect -1181 6 -1177 10
rect -1173 6 -1167 10
rect -1163 6 -1157 10
rect -1153 6 -1147 10
rect -1185 2 -1181 6
rect -1147 2 -1143 6
rect -1171 -6 -1157 2
rect -1084 6 -1080 10
rect -1076 6 -1070 10
rect -1066 6 -1060 10
rect -1056 6 -1050 10
rect -1088 2 -1084 6
rect -1050 2 -1046 6
rect -1074 -6 -1060 2
rect -998 6 -994 10
rect -990 6 -984 10
rect -980 6 -974 10
rect -970 6 -964 10
rect -1002 2 -998 6
rect -964 2 -960 6
rect -988 -6 -974 2
rect -924 6 -920 10
rect -916 6 -910 10
rect -906 6 -900 10
rect -896 6 -890 10
rect -928 2 -924 6
rect -890 2 -886 6
rect -833 8 -829 20
rect -756 10 -752 20
rect -660 10 -656 20
rect -578 10 -574 20
rect -496 10 -492 20
rect -770 6 -766 10
rect -762 6 -756 10
rect -752 6 -746 10
rect -742 6 -736 10
rect -914 -6 -900 2
rect -1265 -22 -1252 -18
rect -1240 -22 -1217 -18
rect -1201 -18 -1183 -14
rect -1240 -28 -1236 -22
rect -1252 -38 -1248 -33
rect -1201 -36 -1197 -18
rect -1166 -21 -1163 -6
rect -1125 -14 -1121 -10
rect -1145 -18 -1121 -14
rect -1100 -18 -1086 -14
rect -1069 -21 -1066 -6
rect -1028 -14 -1024 -10
rect -1048 -18 -1024 -14
rect -1017 -18 -1000 -14
rect -1017 -21 -1014 -18
rect -983 -21 -980 -6
rect -950 -14 -946 -10
rect -962 -18 -946 -14
rect -938 -18 -926 -14
rect -938 -21 -935 -18
rect -909 -21 -906 -6
rect -888 -18 -878 -14
rect -1186 -24 -1118 -21
rect -1186 -27 -1182 -24
rect -1089 -24 -1014 -21
rect -1003 -24 -935 -21
rect -929 -24 -878 -21
rect -1089 -27 -1085 -24
rect -1003 -27 -999 -24
rect -929 -27 -925 -24
rect -1170 -32 -1158 -27
rect -1073 -32 -1061 -27
rect -987 -32 -975 -27
rect -913 -32 -901 -27
rect -881 -28 -878 -24
rect -869 -28 -864 -1
rect -774 2 -770 6
rect -736 2 -732 6
rect -760 -6 -746 2
rect -674 6 -670 10
rect -666 6 -660 10
rect -656 6 -650 10
rect -646 6 -640 10
rect -678 2 -674 6
rect -640 2 -636 6
rect -664 -6 -650 2
rect -592 6 -588 10
rect -584 6 -578 10
rect -574 6 -568 10
rect -564 6 -558 10
rect -596 2 -592 6
rect -558 2 -554 6
rect -582 -6 -568 2
rect -510 6 -506 10
rect -502 6 -496 10
rect -492 6 -486 10
rect -482 6 -476 10
rect -514 2 -510 6
rect -476 2 -472 6
rect -500 -6 -486 2
rect -790 -18 -772 -14
rect -790 -28 -786 -18
rect -755 -21 -752 -6
rect -714 -14 -710 -10
rect -734 -18 -710 -14
rect -690 -18 -676 -14
rect -659 -21 -656 -6
rect -618 -14 -614 -10
rect -638 -18 -614 -14
rect -605 -18 -594 -14
rect -605 -21 -602 -18
rect -577 -21 -574 -6
rect -536 -14 -532 -10
rect -556 -18 -532 -14
rect -525 -18 -512 -14
rect -525 -21 -522 -18
rect -495 -21 -492 -6
rect -474 -18 -464 -14
rect -881 -31 -786 -28
rect -1146 -37 -1142 -32
rect -1252 -45 -1248 -42
rect -1146 -45 -1142 -41
rect -1049 -37 -1045 -32
rect -1049 -45 -1045 -41
rect -963 -37 -959 -32
rect -963 -45 -959 -41
rect -889 -37 -885 -32
rect -790 -36 -786 -31
rect -775 -24 -706 -21
rect -775 -27 -771 -24
rect -679 -24 -602 -21
rect -597 -24 -522 -21
rect -515 -24 -464 -21
rect -679 -27 -675 -24
rect -597 -27 -593 -24
rect -515 -27 -511 -24
rect -759 -32 -747 -27
rect -663 -32 -651 -27
rect -581 -32 -569 -27
rect -499 -32 -487 -27
rect -467 -28 -464 -24
rect -455 -27 -450 -1
rect -455 -28 -409 -27
rect -467 -31 -409 -28
rect -735 -37 -731 -32
rect -889 -45 -885 -41
rect -735 -45 -731 -41
rect -639 -37 -635 -32
rect -639 -45 -635 -41
rect -557 -37 -553 -32
rect -557 -45 -553 -41
rect -475 -37 -471 -32
rect -475 -45 -471 -41
rect -1317 -48 -471 -45
rect -1317 -59 -1287 -54
rect -1234 -123 -1230 -48
rect -1148 -55 -1104 -51
rect -1213 -96 -1209 -65
rect -1196 -73 -1182 -69
rect -1178 -73 -1167 -69
rect -1182 -78 -1178 -73
rect -1170 -96 -1166 -86
rect -1148 -96 -1145 -55
rect -1213 -100 -1182 -96
rect -1170 -100 -1145 -96
rect -1170 -106 -1166 -100
rect -1182 -116 -1178 -111
rect -1182 -123 -1178 -120
rect -823 -119 -819 -48
rect -731 -55 -694 -51
rect -802 -92 -798 -59
rect -785 -69 -771 -65
rect -767 -69 -756 -65
rect -771 -74 -767 -69
rect -759 -92 -755 -82
rect -731 -92 -727 -55
rect -802 -96 -771 -92
rect -759 -96 -727 -92
rect -759 -102 -755 -96
rect -771 -112 -767 -107
rect -771 -119 -767 -116
rect -823 -122 -767 -119
rect -1234 -126 -1178 -123
<< metal2 >>
rect -1310 27 -614 30
rect -1300 -69 -1296 4
rect -1270 -18 -1265 27
rect -1221 20 -1024 23
rect -1221 15 -1217 20
rect -1125 -6 -1121 20
rect -1028 -6 -1024 20
rect -950 20 -864 23
rect -950 -6 -946 20
rect -869 4 -864 20
rect -874 -18 -845 -14
rect -1213 -40 -1201 -36
rect -1213 -54 -1209 -40
rect -1282 -59 -1209 -54
rect -1213 -61 -1209 -59
rect -1118 -65 -1114 -25
rect -1104 -51 -1100 -18
rect -851 -65 -845 -18
rect -1118 -69 -845 -65
rect -833 -65 -829 4
rect -714 -6 -710 27
rect -618 -6 -614 27
rect -536 20 -450 23
rect -536 -6 -532 20
rect -455 4 -450 20
rect -460 -18 -436 -14
rect -802 -40 -790 -36
rect -802 -55 -798 -40
rect -706 -62 -702 -25
rect -694 -51 -690 -18
rect -442 -62 -436 -18
rect -833 -69 -789 -65
rect -706 -66 -436 -62
rect -1300 -73 -1200 -69
<< ntransistor >>
rect -1245 -33 -1243 -29
rect -1179 -31 -1177 -27
rect -1151 -31 -1149 -27
rect -1082 -31 -1080 -27
rect -1054 -31 -1052 -27
rect -996 -31 -994 -27
rect -968 -31 -966 -27
rect -922 -31 -920 -27
rect -894 -31 -892 -27
rect -768 -31 -766 -27
rect -740 -31 -738 -27
rect -672 -31 -670 -27
rect -644 -31 -642 -27
rect -590 -31 -588 -27
rect -562 -31 -560 -27
rect -508 -31 -506 -27
rect -480 -31 -478 -27
rect -1175 -111 -1173 -107
rect -764 -107 -762 -103
<< ptransistor >>
rect -1245 -8 -1243 0
rect -1179 -6 -1177 2
rect -1151 -6 -1149 2
rect -1082 -6 -1080 2
rect -1054 -6 -1052 2
rect -996 -6 -994 2
rect -968 -6 -966 2
rect -922 -6 -920 2
rect -894 -6 -892 2
rect -768 -6 -766 2
rect -740 -6 -738 2
rect -672 -6 -670 2
rect -644 -6 -642 2
rect -590 -6 -588 2
rect -562 -6 -560 2
rect -508 -6 -506 2
rect -480 -6 -478 2
rect -1175 -86 -1173 -78
rect -764 -82 -762 -74
<< polycontact >>
rect -1252 -22 -1248 -18
rect -1183 -18 -1179 -14
rect -1149 -18 -1145 -14
rect -1086 -18 -1082 -14
rect -1052 -18 -1048 -14
rect -1000 -18 -996 -14
rect -966 -18 -962 -14
rect -926 -18 -922 -14
rect -892 -18 -888 -14
rect -772 -18 -768 -14
rect -738 -18 -734 -14
rect -676 -18 -672 -14
rect -642 -18 -638 -14
rect -594 -18 -590 -14
rect -560 -18 -556 -14
rect -512 -18 -508 -14
rect -478 -18 -474 -14
rect -1182 -100 -1178 -96
rect -771 -96 -767 -92
<< ndcontact >>
rect -1252 -33 -1248 -28
rect -1240 -33 -1236 -28
rect -1186 -32 -1182 -27
rect -1174 -32 -1170 -27
rect -1158 -32 -1154 -27
rect -1146 -32 -1142 -27
rect -1089 -32 -1085 -27
rect -1077 -32 -1073 -27
rect -1061 -32 -1057 -27
rect -1049 -32 -1045 -27
rect -1003 -32 -999 -27
rect -991 -32 -987 -27
rect -975 -32 -971 -27
rect -963 -32 -959 -27
rect -929 -32 -925 -27
rect -917 -32 -913 -27
rect -901 -32 -897 -27
rect -889 -32 -885 -27
rect -775 -32 -771 -27
rect -763 -32 -759 -27
rect -747 -32 -743 -27
rect -735 -32 -731 -27
rect -679 -32 -675 -27
rect -667 -32 -663 -27
rect -651 -32 -647 -27
rect -639 -32 -635 -27
rect -597 -32 -593 -27
rect -585 -32 -581 -27
rect -569 -32 -565 -27
rect -557 -32 -553 -27
rect -515 -32 -511 -27
rect -503 -32 -499 -27
rect -487 -32 -483 -27
rect -475 -32 -471 -27
rect -1182 -111 -1178 -106
rect -1170 -111 -1166 -106
rect -771 -107 -767 -102
rect -759 -107 -755 -102
<< pdcontact >>
rect -1252 -8 -1248 0
rect -1240 -8 -1236 0
rect -1185 -6 -1181 2
rect -1175 -6 -1171 2
rect -1157 -6 -1153 2
rect -1147 -6 -1143 2
rect -1088 -6 -1084 2
rect -1078 -6 -1074 2
rect -1060 -6 -1056 2
rect -1050 -6 -1046 2
rect -1002 -6 -998 2
rect -992 -6 -988 2
rect -974 -6 -970 2
rect -964 -6 -960 2
rect -928 -6 -924 2
rect -918 -6 -914 2
rect -900 -6 -896 2
rect -890 -6 -886 2
rect -774 -6 -770 2
rect -764 -6 -760 2
rect -746 -6 -742 2
rect -736 -6 -732 2
rect -678 -6 -674 2
rect -668 -6 -664 2
rect -650 -6 -646 2
rect -640 -6 -636 2
rect -596 -6 -592 2
rect -586 -6 -582 2
rect -568 -6 -564 2
rect -558 -6 -554 2
rect -514 -6 -510 2
rect -504 -6 -500 2
rect -486 -6 -482 2
rect -476 -6 -472 2
rect -1182 -86 -1178 -78
rect -1170 -86 -1166 -78
rect -771 -82 -767 -74
rect -759 -82 -755 -74
<< m2contact >>
rect -1300 4 -1296 8
rect -1221 11 -1217 15
rect -833 4 -829 8
rect -869 -1 -864 4
rect -1270 -22 -1265 -18
rect -1125 -10 -1121 -6
rect -1104 -18 -1100 -14
rect -1028 -10 -1024 -6
rect -950 -10 -946 -6
rect -878 -18 -874 -14
rect -1118 -25 -1114 -21
rect -455 -1 -450 4
rect -714 -10 -710 -6
rect -694 -18 -690 -14
rect -618 -10 -614 -6
rect -536 -10 -532 -6
rect -464 -18 -460 -14
rect -1201 -40 -1197 -36
rect -706 -25 -702 -21
rect -790 -40 -786 -36
rect -1287 -59 -1282 -54
rect -1104 -55 -1100 -51
rect -1213 -65 -1209 -61
rect -1200 -73 -1196 -69
rect -694 -55 -690 -51
rect -802 -59 -798 -55
rect -789 -69 -785 -65
<< psubstratepcontact >>
rect -1252 -42 -1248 -38
rect -1146 -41 -1142 -37
rect -1049 -41 -1045 -37
rect -963 -41 -959 -37
rect -889 -41 -885 -37
rect -735 -41 -731 -37
rect -639 -41 -635 -37
rect -557 -41 -553 -37
rect -475 -41 -471 -37
rect -771 -116 -767 -112
rect -1182 -120 -1178 -116
<< nsubstratencontact >>
rect -1252 5 -1248 9
rect -1237 5 -1233 9
rect -1185 6 -1181 10
rect -1177 6 -1173 10
rect -1167 6 -1163 10
rect -1157 6 -1153 10
rect -1147 6 -1143 10
rect -1088 6 -1084 10
rect -1080 6 -1076 10
rect -1070 6 -1066 10
rect -1060 6 -1056 10
rect -1050 6 -1046 10
rect -1002 6 -998 10
rect -994 6 -990 10
rect -984 6 -980 10
rect -974 6 -970 10
rect -964 6 -960 10
rect -928 6 -924 10
rect -920 6 -916 10
rect -910 6 -906 10
rect -900 6 -896 10
rect -890 6 -886 10
rect -774 6 -770 10
rect -766 6 -762 10
rect -756 6 -752 10
rect -746 6 -742 10
rect -736 6 -732 10
rect -678 6 -674 10
rect -670 6 -666 10
rect -660 6 -656 10
rect -650 6 -646 10
rect -640 6 -636 10
rect -596 6 -592 10
rect -588 6 -584 10
rect -578 6 -574 10
rect -568 6 -564 10
rect -558 6 -554 10
rect -514 6 -510 10
rect -506 6 -502 10
rect -496 6 -492 10
rect -486 6 -482 10
rect -476 6 -472 10
rect -771 -69 -767 -65
rect -756 -69 -752 -65
rect -1182 -73 -1178 -69
rect -1167 -73 -1163 -69
<< labels >>
rlabel m2contact -1221 15 -1217 15 1 invout
rlabel metal1 -1236 -22 -1236 -17 1 invout
rlabel pdcontact -1185 1 -1185 1 1 M6source
rlabel pdcontact -1145 0 -1145 0 1 M7source
rlabel pdcontact -1088 1 -1088 1 1 M6source
rlabel pdcontact -1048 0 -1048 0 1 M7source
rlabel pdcontact -1002 1 -1002 1 1 M6source
rlabel pdcontact -962 0 -962 0 1 M7source
rlabel pdcontact -928 1 -928 1 1 M6source
rlabel pdcontact -888 0 -888 0 1 M7source
rlabel pdcontact -774 1 -774 1 1 M6source
rlabel pdcontact -734 0 -734 0 1 M7source
rlabel pdcontact -678 1 -678 1 1 M6source
rlabel pdcontact -638 0 -638 0 1 M7source
rlabel pdcontact -596 1 -596 1 1 M6source
rlabel pdcontact -556 0 -556 0 1 M7source
rlabel pdcontact -514 1 -514 1 1 M6source
rlabel pdcontact -474 0 -474 0 1 M7source
rlabel metal1 -1317 -48 -1317 -45 3 gnd!
rlabel metal1 -1317 -59 -1317 -54 3 D
rlabel metal1 -1311 20 -1311 23 1 vdd!
rlabel metal2 -1310 27 -1310 30 5 clock
rlabel metal1 -409 -31 -409 -27 7 out
<< end >>
