magic
tech scmos
timestamp 1398365948
<< nwell >>
rect -66 -10 -38 15
rect 2 -7 55 18
rect 138 -7 191 18
rect 303 -7 356 18
rect 444 -7 497 18
rect 4 -101 32 -76
<< polysilicon >>
rect 13 7 15 9
rect 41 7 43 9
rect 149 7 151 9
rect 177 7 179 9
rect 314 7 316 9
rect 342 7 344 9
rect 455 7 457 9
rect 483 7 485 9
rect -53 5 -51 7
rect -53 -14 -51 -3
rect -56 -16 -51 -14
rect -53 -24 -51 -16
rect 13 -22 15 -1
rect 41 -22 43 -1
rect 149 -22 151 -1
rect 177 -22 179 -1
rect 314 -22 316 -1
rect 342 -22 344 -1
rect 455 -22 457 -1
rect 483 -22 485 -1
rect 13 -28 15 -26
rect 41 -28 43 -26
rect 149 -28 151 -26
rect 177 -28 179 -26
rect 314 -28 316 -26
rect 342 -28 344 -26
rect 455 -28 457 -26
rect 483 -28 485 -26
rect -53 -30 -51 -28
rect 17 -86 19 -84
rect 17 -105 19 -94
rect 14 -107 19 -105
rect 17 -115 19 -107
rect 17 -121 19 -119
<< ndiffusion >>
rect -56 -28 -53 -24
rect -51 -28 -48 -24
rect 10 -26 13 -22
rect 15 -26 18 -22
rect 38 -26 41 -22
rect 43 -26 46 -22
rect 146 -26 149 -22
rect 151 -26 154 -22
rect 174 -26 177 -22
rect 179 -26 182 -22
rect 311 -26 314 -22
rect 316 -26 319 -22
rect 339 -26 342 -22
rect 344 -26 347 -22
rect 452 -26 455 -22
rect 457 -26 460 -22
rect 480 -26 483 -22
rect 485 -26 488 -22
rect 14 -119 17 -115
rect 19 -119 22 -115
<< pdiffusion >>
rect -56 -3 -53 5
rect -51 -3 -48 5
rect 11 -1 13 7
rect 15 -1 17 7
rect 39 -1 41 7
rect 43 -1 45 7
rect 147 -1 149 7
rect 151 -1 153 7
rect 175 -1 177 7
rect 179 -1 181 7
rect 312 -1 314 7
rect 316 -1 318 7
rect 340 -1 342 7
rect 344 -1 346 7
rect 453 -1 455 7
rect 457 -1 459 7
rect 481 -1 483 7
rect 485 -1 487 7
rect 14 -94 17 -86
rect 19 -94 22 -86
<< metal1 >>
rect -135 25 471 28
rect -108 13 -104 25
rect -45 14 -41 25
rect -56 10 -45 14
rect -60 5 -56 10
rect -48 -13 -44 -3
rect -29 -13 -25 16
rect 25 15 29 25
rect 161 15 165 25
rect 326 15 330 21
rect 467 15 471 25
rect 11 11 15 15
rect 19 11 25 15
rect 29 11 35 15
rect 39 11 45 15
rect 7 7 11 11
rect 45 7 49 11
rect 21 -1 35 7
rect 147 11 151 15
rect 155 11 161 15
rect 165 11 171 15
rect 175 11 181 15
rect 143 7 147 11
rect 181 7 185 11
rect 157 -1 171 7
rect 312 11 316 15
rect 320 11 326 15
rect 330 11 336 15
rect 340 11 346 15
rect 308 7 312 11
rect 346 7 350 11
rect 322 -1 336 7
rect 453 11 457 15
rect 461 11 467 15
rect 471 11 477 15
rect 481 11 487 15
rect 449 7 453 11
rect 487 7 491 11
rect 463 -1 477 7
rect -76 -17 -60 -13
rect -48 -17 -25 -13
rect -9 -13 9 -9
rect -48 -23 -44 -17
rect -60 -33 -56 -28
rect -9 -31 -5 -13
rect 26 -16 29 -1
rect 67 -9 71 -5
rect 47 -13 71 -9
rect 119 -13 145 -9
rect 162 -16 165 -1
rect 203 -9 207 -5
rect 183 -13 207 -9
rect 293 -13 310 -9
rect 293 -16 296 -13
rect 327 -16 330 -1
rect 368 -9 372 -5
rect 348 -13 372 -9
rect 430 -13 451 -9
rect 430 -16 433 -13
rect 468 -16 471 -1
rect 489 -13 499 -9
rect 6 -19 87 -16
rect 6 -22 10 -19
rect 142 -19 296 -16
rect 307 -19 433 -16
rect 448 -19 499 -16
rect 142 -22 146 -19
rect 307 -22 311 -19
rect 448 -22 452 -19
rect 22 -27 34 -22
rect 158 -27 170 -22
rect 323 -27 335 -22
rect 464 -27 476 -22
rect 496 -23 499 -19
rect 508 -23 513 4
rect 496 -26 521 -23
rect 46 -32 50 -27
rect -60 -40 -56 -37
rect 46 -40 50 -36
rect 182 -32 186 -27
rect 182 -40 186 -36
rect 347 -32 351 -27
rect 347 -40 351 -36
rect 488 -32 492 -27
rect 488 -40 492 -36
rect -122 -43 492 -40
rect -129 -54 -95 -49
rect -42 -131 -38 -43
rect -21 -104 -17 -64
rect -4 -81 10 -77
rect 14 -81 25 -77
rect 10 -86 14 -81
rect 22 -104 26 -94
rect 115 -104 119 -60
rect -21 -108 10 -104
rect 22 -108 119 -104
rect 22 -114 26 -108
rect 10 -124 14 -119
rect 10 -131 14 -128
rect -42 -134 14 -131
<< metal2 >>
rect -29 38 207 41
rect -29 20 -25 38
rect -108 -77 -104 9
rect 67 -1 71 38
rect 203 -1 207 38
rect 368 36 513 40
rect 368 -1 372 36
rect 508 9 513 36
rect 503 -13 545 -9
rect -21 -35 -9 -31
rect -21 -49 -17 -35
rect -90 -54 -17 -49
rect -21 -60 -17 -54
rect 87 -74 91 -20
rect 115 -56 119 -13
rect 539 -74 545 -13
rect 87 -77 545 -74
rect -108 -81 -8 -77
rect 88 -78 545 -77
<< ntransistor >>
rect -53 -28 -51 -24
rect 13 -26 15 -22
rect 41 -26 43 -22
rect 149 -26 151 -22
rect 177 -26 179 -22
rect 314 -26 316 -22
rect 342 -26 344 -22
rect 455 -26 457 -22
rect 483 -26 485 -22
rect 17 -119 19 -115
<< ptransistor >>
rect -53 -3 -51 5
rect 13 -1 15 7
rect 41 -1 43 7
rect 149 -1 151 7
rect 177 -1 179 7
rect 314 -1 316 7
rect 342 -1 344 7
rect 455 -1 457 7
rect 483 -1 485 7
rect 17 -94 19 -86
<< polycontact >>
rect -60 -17 -56 -13
rect 9 -13 13 -9
rect 43 -13 47 -9
rect 145 -13 149 -9
rect 179 -13 183 -9
rect 310 -13 314 -9
rect 344 -13 348 -9
rect 451 -13 455 -9
rect 485 -13 489 -9
rect 10 -108 14 -104
<< ndcontact >>
rect -60 -28 -56 -23
rect -48 -28 -44 -23
rect 6 -27 10 -22
rect 18 -27 22 -22
rect 34 -27 38 -22
rect 46 -27 50 -22
rect 142 -27 146 -22
rect 154 -27 158 -22
rect 170 -27 174 -22
rect 182 -27 186 -22
rect 307 -27 311 -22
rect 319 -27 323 -22
rect 335 -27 339 -22
rect 347 -27 351 -22
rect 448 -27 452 -22
rect 460 -27 464 -22
rect 476 -27 480 -22
rect 488 -27 492 -22
rect 10 -119 14 -114
rect 22 -119 26 -114
<< pdcontact >>
rect -60 -3 -56 5
rect -48 -3 -44 5
rect 7 -1 11 7
rect 17 -1 21 7
rect 35 -1 39 7
rect 45 -1 49 7
rect 143 -1 147 7
rect 153 -1 157 7
rect 171 -1 175 7
rect 181 -1 185 7
rect 308 -1 312 7
rect 318 -1 322 7
rect 336 -1 340 7
rect 346 -1 350 7
rect 449 -1 453 7
rect 459 -1 463 7
rect 477 -1 481 7
rect 487 -1 491 7
rect 10 -94 14 -86
rect 22 -94 26 -86
<< m2contact >>
rect -108 9 -104 13
rect -29 16 -25 20
rect 508 4 513 9
rect 67 -5 71 -1
rect 115 -13 119 -9
rect 203 -5 207 -1
rect 368 -5 372 -1
rect 499 -13 503 -9
rect 87 -20 91 -16
rect -9 -35 -5 -31
rect -95 -54 -90 -49
rect 115 -60 119 -56
rect -21 -64 -17 -60
rect -8 -81 -4 -77
<< psubstratepcontact >>
rect -60 -37 -56 -33
rect 46 -36 50 -32
rect 182 -36 186 -32
rect 347 -36 351 -32
rect 488 -36 492 -32
rect 10 -128 14 -124
<< nsubstratencontact >>
rect -60 10 -56 14
rect -45 10 -41 14
rect 7 11 11 15
rect 15 11 19 15
rect 25 11 29 15
rect 35 11 39 15
rect 45 11 49 15
rect 143 11 147 15
rect 151 11 155 15
rect 161 11 165 15
rect 171 11 175 15
rect 181 11 185 15
rect 308 11 312 15
rect 316 11 320 15
rect 326 11 330 15
rect 336 11 340 15
rect 346 11 350 15
rect 449 11 453 15
rect 457 11 461 15
rect 467 11 471 15
rect 477 11 481 15
rect 487 11 491 15
rect 10 -81 14 -77
rect 25 -81 29 -77
<< labels >>
rlabel metal1 -76 -17 -76 -13 1 clock
rlabel m2contact -29 20 -25 20 1 invout
rlabel metal1 -44 -17 -44 -12 1 invout
rlabel pdcontact 7 6 7 6 1 M6source
rlabel pdcontact 47 5 47 5 1 M7source
rlabel pdcontact 143 6 143 6 1 M6source
rlabel pdcontact 183 5 183 5 1 M7source
rlabel metal1 -135 25 -135 28 3 vdd!
rlabel metal1 -122 -43 -122 -40 1 gnd!
rlabel pdcontact 449 6 449 6 1 M6source
rlabel pdcontact 489 5 489 5 1 M7source
rlabel pdcontact 308 6 308 6 1 M6source
rlabel pdcontact 348 5 348 5 1 M7source
rlabel metal1 521 -26 521 -23 7 Q
rlabel metal1 -129 -54 -129 -49 1 D
<< end >>
