magic
tech scmos
timestamp 1398872030
<< nwell >>
rect -1244 24 -1216 49
rect -1176 27 -1123 52
rect -1079 27 -1026 52
rect -993 27 -940 52
rect -919 27 -866 52
rect -765 27 -712 52
rect -669 27 -616 52
rect -587 27 -534 52
rect -505 27 -452 52
rect -1174 -54 -1146 -29
rect -763 -50 -735 -25
rect -1244 -168 -1216 -143
rect -1176 -165 -1123 -140
rect -1079 -165 -1026 -140
rect -993 -165 -940 -140
rect -919 -165 -866 -140
rect -765 -165 -712 -140
rect -669 -165 -616 -140
rect -587 -165 -534 -140
rect -505 -165 -452 -140
rect -1174 -246 -1146 -221
rect -763 -242 -735 -217
rect -1244 -359 -1216 -334
rect -1176 -356 -1123 -331
rect -1079 -356 -1026 -331
rect -993 -356 -940 -331
rect -919 -356 -866 -331
rect -765 -356 -712 -331
rect -669 -356 -616 -331
rect -587 -356 -534 -331
rect -505 -356 -452 -331
rect -1174 -437 -1146 -412
rect -763 -433 -735 -408
rect -1245 -545 -1217 -520
rect -1177 -542 -1124 -517
rect -1080 -542 -1027 -517
rect -994 -542 -941 -517
rect -920 -542 -867 -517
rect -766 -542 -713 -517
rect -670 -542 -617 -517
rect -588 -542 -535 -517
rect -506 -542 -453 -517
rect -1175 -623 -1147 -598
rect -764 -619 -736 -594
rect -1227 -715 -1174 -690
rect -1144 -715 -1091 -690
rect -1037 -715 -984 -690
rect -954 -715 -901 -690
<< polysilicon >>
rect -1165 41 -1163 43
rect -1137 41 -1135 43
rect -1068 41 -1066 43
rect -1040 41 -1038 43
rect -982 41 -980 43
rect -954 41 -952 43
rect -908 41 -906 43
rect -880 41 -878 43
rect -754 41 -752 43
rect -726 41 -724 43
rect -658 41 -656 43
rect -630 41 -628 43
rect -576 41 -574 43
rect -548 41 -546 43
rect -494 41 -492 43
rect -466 41 -464 43
rect -1231 39 -1229 41
rect -1231 20 -1229 31
rect -1234 18 -1229 20
rect -1231 10 -1229 18
rect -1165 11 -1163 33
rect -1137 11 -1135 33
rect -1068 11 -1066 33
rect -1040 11 -1038 33
rect -982 11 -980 33
rect -954 11 -952 33
rect -908 11 -906 33
rect -880 11 -878 33
rect -754 11 -752 33
rect -726 11 -724 33
rect -658 12 -656 33
rect -630 12 -628 33
rect -576 11 -574 33
rect -548 11 -546 33
rect -494 11 -492 33
rect -466 11 -464 33
rect -1231 4 -1229 6
rect -1165 5 -1163 7
rect -1137 5 -1135 7
rect -1068 5 -1066 7
rect -1040 5 -1038 7
rect -982 5 -980 7
rect -954 5 -952 7
rect -908 5 -906 7
rect -880 5 -878 7
rect -754 5 -752 7
rect -726 5 -724 7
rect -658 6 -656 8
rect -630 6 -628 8
rect -576 5 -574 7
rect -548 5 -546 7
rect -494 5 -492 7
rect -466 5 -464 7
rect -750 -35 -748 -33
rect -1161 -39 -1159 -37
rect -1161 -58 -1159 -47
rect -750 -54 -748 -43
rect -753 -56 -748 -54
rect -1164 -60 -1159 -58
rect -1161 -68 -1159 -60
rect -750 -64 -748 -56
rect -750 -70 -748 -68
rect -1161 -74 -1159 -72
rect -1165 -151 -1163 -149
rect -1137 -151 -1135 -149
rect -1068 -151 -1066 -149
rect -1040 -151 -1038 -149
rect -982 -151 -980 -149
rect -954 -151 -952 -149
rect -908 -151 -906 -149
rect -880 -151 -878 -149
rect -754 -151 -752 -149
rect -726 -151 -724 -149
rect -658 -151 -656 -149
rect -630 -151 -628 -149
rect -576 -151 -574 -149
rect -548 -151 -546 -149
rect -494 -151 -492 -149
rect -466 -151 -464 -149
rect -1231 -153 -1229 -151
rect -1231 -172 -1229 -161
rect -1234 -174 -1229 -172
rect -1231 -182 -1229 -174
rect -1165 -181 -1163 -159
rect -1137 -181 -1135 -159
rect -1068 -181 -1066 -159
rect -1040 -181 -1038 -159
rect -982 -181 -980 -159
rect -954 -181 -952 -159
rect -908 -181 -906 -159
rect -880 -181 -878 -159
rect -754 -181 -752 -159
rect -726 -181 -724 -159
rect -658 -180 -656 -159
rect -630 -180 -628 -159
rect -576 -181 -574 -159
rect -548 -181 -546 -159
rect -494 -181 -492 -159
rect -466 -181 -464 -159
rect -1231 -188 -1229 -186
rect -1165 -187 -1163 -185
rect -1137 -187 -1135 -185
rect -1068 -187 -1066 -185
rect -1040 -187 -1038 -185
rect -982 -187 -980 -185
rect -954 -187 -952 -185
rect -908 -187 -906 -185
rect -880 -187 -878 -185
rect -754 -187 -752 -185
rect -726 -187 -724 -185
rect -658 -186 -656 -184
rect -630 -186 -628 -184
rect -576 -187 -574 -185
rect -548 -187 -546 -185
rect -494 -187 -492 -185
rect -466 -187 -464 -185
rect -750 -227 -748 -225
rect -1161 -231 -1159 -229
rect -1161 -250 -1159 -239
rect -750 -246 -748 -235
rect -753 -248 -748 -246
rect -1164 -252 -1159 -250
rect -1161 -260 -1159 -252
rect -750 -256 -748 -248
rect -750 -262 -748 -260
rect -1161 -266 -1159 -264
rect -1165 -342 -1163 -340
rect -1137 -342 -1135 -340
rect -1068 -342 -1066 -340
rect -1040 -342 -1038 -340
rect -982 -342 -980 -340
rect -954 -342 -952 -340
rect -908 -342 -906 -340
rect -880 -342 -878 -340
rect -754 -342 -752 -340
rect -726 -342 -724 -340
rect -658 -342 -656 -340
rect -630 -342 -628 -340
rect -576 -342 -574 -340
rect -548 -342 -546 -340
rect -494 -342 -492 -340
rect -466 -342 -464 -340
rect -1231 -344 -1229 -342
rect -1231 -363 -1229 -352
rect -1234 -365 -1229 -363
rect -1231 -373 -1229 -365
rect -1165 -372 -1163 -350
rect -1137 -372 -1135 -350
rect -1068 -372 -1066 -350
rect -1040 -372 -1038 -350
rect -982 -372 -980 -350
rect -954 -372 -952 -350
rect -908 -372 -906 -350
rect -880 -372 -878 -350
rect -754 -372 -752 -350
rect -726 -372 -724 -350
rect -658 -371 -656 -350
rect -630 -371 -628 -350
rect -576 -372 -574 -350
rect -548 -372 -546 -350
rect -494 -372 -492 -350
rect -466 -372 -464 -350
rect -1231 -379 -1229 -377
rect -1165 -378 -1163 -376
rect -1137 -378 -1135 -376
rect -1068 -378 -1066 -376
rect -1040 -378 -1038 -376
rect -982 -378 -980 -376
rect -954 -378 -952 -376
rect -908 -378 -906 -376
rect -880 -378 -878 -376
rect -754 -378 -752 -376
rect -726 -378 -724 -376
rect -658 -377 -656 -375
rect -630 -377 -628 -375
rect -576 -378 -574 -376
rect -548 -378 -546 -376
rect -494 -378 -492 -376
rect -466 -378 -464 -376
rect -750 -418 -748 -416
rect -1161 -422 -1159 -420
rect -1161 -441 -1159 -430
rect -750 -437 -748 -426
rect -753 -439 -748 -437
rect -1164 -443 -1159 -441
rect -1161 -451 -1159 -443
rect -750 -447 -748 -439
rect -750 -453 -748 -451
rect -1161 -457 -1159 -455
rect -1166 -528 -1164 -526
rect -1138 -528 -1136 -526
rect -1069 -528 -1067 -526
rect -1041 -528 -1039 -526
rect -983 -528 -981 -526
rect -955 -528 -953 -526
rect -909 -528 -907 -526
rect -881 -528 -879 -526
rect -755 -528 -753 -526
rect -727 -528 -725 -526
rect -659 -528 -657 -526
rect -631 -528 -629 -526
rect -577 -528 -575 -526
rect -549 -528 -547 -526
rect -495 -528 -493 -526
rect -467 -528 -465 -526
rect -1232 -530 -1230 -528
rect -1232 -549 -1230 -538
rect -1235 -551 -1230 -549
rect -1232 -559 -1230 -551
rect -1166 -558 -1164 -536
rect -1138 -558 -1136 -536
rect -1069 -558 -1067 -536
rect -1041 -558 -1039 -536
rect -983 -558 -981 -536
rect -955 -558 -953 -536
rect -909 -558 -907 -536
rect -881 -558 -879 -536
rect -755 -558 -753 -536
rect -727 -558 -725 -536
rect -659 -557 -657 -536
rect -631 -557 -629 -536
rect -577 -558 -575 -536
rect -549 -558 -547 -536
rect -495 -558 -493 -536
rect -467 -558 -465 -536
rect -1232 -565 -1230 -563
rect -1166 -564 -1164 -562
rect -1138 -564 -1136 -562
rect -1069 -564 -1067 -562
rect -1041 -564 -1039 -562
rect -983 -564 -981 -562
rect -955 -564 -953 -562
rect -909 -564 -907 -562
rect -881 -564 -879 -562
rect -755 -564 -753 -562
rect -727 -564 -725 -562
rect -659 -563 -657 -561
rect -631 -563 -629 -561
rect -577 -564 -575 -562
rect -549 -564 -547 -562
rect -495 -564 -493 -562
rect -467 -564 -465 -562
rect -751 -604 -749 -602
rect -1162 -608 -1160 -606
rect -1162 -627 -1160 -616
rect -751 -623 -749 -612
rect -754 -625 -749 -623
rect -1165 -629 -1160 -627
rect -1162 -637 -1160 -629
rect -751 -633 -749 -625
rect -751 -639 -749 -637
rect -1162 -643 -1160 -641
rect -1216 -701 -1214 -699
rect -1188 -701 -1186 -699
rect -1133 -701 -1131 -699
rect -1105 -701 -1103 -699
rect -1026 -701 -1024 -699
rect -998 -701 -996 -699
rect -943 -701 -941 -699
rect -915 -701 -913 -699
rect -1216 -731 -1214 -709
rect -1188 -731 -1186 -709
rect -1133 -731 -1131 -709
rect -1105 -731 -1103 -709
rect -1026 -731 -1024 -709
rect -998 -731 -996 -709
rect -943 -731 -941 -709
rect -915 -731 -913 -709
rect -1216 -737 -1214 -735
rect -1188 -737 -1186 -735
rect -1133 -737 -1131 -735
rect -1105 -737 -1103 -735
rect -1026 -737 -1024 -735
rect -998 -737 -996 -735
rect -943 -737 -941 -735
rect -915 -737 -913 -735
<< ndiffusion >>
rect -1234 6 -1231 10
rect -1229 6 -1226 10
rect -1168 7 -1165 11
rect -1163 7 -1160 11
rect -1140 7 -1137 11
rect -1135 7 -1132 11
rect -1071 7 -1068 11
rect -1066 7 -1063 11
rect -1043 7 -1040 11
rect -1038 7 -1035 11
rect -985 7 -982 11
rect -980 7 -977 11
rect -957 7 -954 11
rect -952 7 -949 11
rect -911 7 -908 11
rect -906 7 -903 11
rect -883 7 -880 11
rect -878 7 -875 11
rect -757 7 -754 11
rect -752 7 -749 11
rect -729 7 -726 11
rect -724 7 -721 11
rect -661 8 -658 12
rect -656 8 -653 12
rect -633 8 -630 12
rect -628 8 -625 12
rect -579 7 -576 11
rect -574 7 -571 11
rect -551 7 -548 11
rect -546 7 -543 11
rect -497 7 -494 11
rect -492 7 -489 11
rect -469 7 -466 11
rect -464 7 -461 11
rect -753 -68 -750 -64
rect -748 -68 -745 -64
rect -1164 -72 -1161 -68
rect -1159 -72 -1156 -68
rect -1234 -186 -1231 -182
rect -1229 -186 -1226 -182
rect -1168 -185 -1165 -181
rect -1163 -185 -1160 -181
rect -1140 -185 -1137 -181
rect -1135 -185 -1132 -181
rect -1071 -185 -1068 -181
rect -1066 -185 -1063 -181
rect -1043 -185 -1040 -181
rect -1038 -185 -1035 -181
rect -985 -185 -982 -181
rect -980 -185 -977 -181
rect -957 -185 -954 -181
rect -952 -185 -949 -181
rect -911 -185 -908 -181
rect -906 -185 -903 -181
rect -883 -185 -880 -181
rect -878 -185 -875 -181
rect -757 -185 -754 -181
rect -752 -185 -749 -181
rect -729 -185 -726 -181
rect -724 -185 -721 -181
rect -661 -184 -658 -180
rect -656 -184 -653 -180
rect -633 -184 -630 -180
rect -628 -184 -625 -180
rect -579 -185 -576 -181
rect -574 -185 -571 -181
rect -551 -185 -548 -181
rect -546 -185 -543 -181
rect -497 -185 -494 -181
rect -492 -185 -489 -181
rect -469 -185 -466 -181
rect -464 -185 -461 -181
rect -753 -260 -750 -256
rect -748 -260 -745 -256
rect -1164 -264 -1161 -260
rect -1159 -264 -1156 -260
rect -1234 -377 -1231 -373
rect -1229 -377 -1226 -373
rect -1168 -376 -1165 -372
rect -1163 -376 -1160 -372
rect -1140 -376 -1137 -372
rect -1135 -376 -1132 -372
rect -1071 -376 -1068 -372
rect -1066 -376 -1063 -372
rect -1043 -376 -1040 -372
rect -1038 -376 -1035 -372
rect -985 -376 -982 -372
rect -980 -376 -977 -372
rect -957 -376 -954 -372
rect -952 -376 -949 -372
rect -911 -376 -908 -372
rect -906 -376 -903 -372
rect -883 -376 -880 -372
rect -878 -376 -875 -372
rect -757 -376 -754 -372
rect -752 -376 -749 -372
rect -729 -376 -726 -372
rect -724 -376 -721 -372
rect -661 -375 -658 -371
rect -656 -375 -653 -371
rect -633 -375 -630 -371
rect -628 -375 -625 -371
rect -579 -376 -576 -372
rect -574 -376 -571 -372
rect -551 -376 -548 -372
rect -546 -376 -543 -372
rect -497 -376 -494 -372
rect -492 -376 -489 -372
rect -469 -376 -466 -372
rect -464 -376 -461 -372
rect -753 -451 -750 -447
rect -748 -451 -745 -447
rect -1164 -455 -1161 -451
rect -1159 -455 -1156 -451
rect -1235 -563 -1232 -559
rect -1230 -563 -1227 -559
rect -1169 -562 -1166 -558
rect -1164 -562 -1161 -558
rect -1141 -562 -1138 -558
rect -1136 -562 -1133 -558
rect -1072 -562 -1069 -558
rect -1067 -562 -1064 -558
rect -1044 -562 -1041 -558
rect -1039 -562 -1036 -558
rect -986 -562 -983 -558
rect -981 -562 -978 -558
rect -958 -562 -955 -558
rect -953 -562 -950 -558
rect -912 -562 -909 -558
rect -907 -562 -904 -558
rect -884 -562 -881 -558
rect -879 -562 -876 -558
rect -758 -562 -755 -558
rect -753 -562 -750 -558
rect -730 -562 -727 -558
rect -725 -562 -722 -558
rect -662 -561 -659 -557
rect -657 -561 -654 -557
rect -634 -561 -631 -557
rect -629 -561 -626 -557
rect -580 -562 -577 -558
rect -575 -562 -572 -558
rect -552 -562 -549 -558
rect -547 -562 -544 -558
rect -498 -562 -495 -558
rect -493 -562 -490 -558
rect -470 -562 -467 -558
rect -465 -562 -462 -558
rect -754 -637 -751 -633
rect -749 -637 -746 -633
rect -1165 -641 -1162 -637
rect -1160 -641 -1157 -637
rect -1219 -735 -1216 -731
rect -1214 -735 -1211 -731
rect -1191 -735 -1188 -731
rect -1186 -735 -1183 -731
rect -1136 -735 -1133 -731
rect -1131 -735 -1128 -731
rect -1108 -735 -1105 -731
rect -1103 -735 -1100 -731
rect -1029 -735 -1026 -731
rect -1024 -735 -1021 -731
rect -1001 -735 -998 -731
rect -996 -735 -993 -731
rect -946 -735 -943 -731
rect -941 -735 -938 -731
rect -918 -735 -915 -731
rect -913 -735 -910 -731
<< pdiffusion >>
rect -1234 31 -1231 39
rect -1229 31 -1226 39
rect -1167 33 -1165 41
rect -1163 33 -1161 41
rect -1139 33 -1137 41
rect -1135 33 -1133 41
rect -1070 33 -1068 41
rect -1066 33 -1064 41
rect -1042 33 -1040 41
rect -1038 33 -1036 41
rect -984 33 -982 41
rect -980 33 -978 41
rect -956 33 -954 41
rect -952 33 -950 41
rect -910 33 -908 41
rect -906 33 -904 41
rect -882 33 -880 41
rect -878 33 -876 41
rect -756 33 -754 41
rect -752 33 -750 41
rect -728 33 -726 41
rect -724 33 -722 41
rect -660 33 -658 41
rect -656 33 -654 41
rect -632 33 -630 41
rect -628 33 -626 41
rect -578 33 -576 41
rect -574 33 -572 41
rect -550 33 -548 41
rect -546 33 -544 41
rect -496 33 -494 41
rect -492 33 -490 41
rect -468 33 -466 41
rect -464 33 -462 41
rect -1164 -47 -1161 -39
rect -1159 -47 -1156 -39
rect -753 -43 -750 -35
rect -748 -43 -745 -35
rect -1234 -161 -1231 -153
rect -1229 -161 -1226 -153
rect -1167 -159 -1165 -151
rect -1163 -159 -1161 -151
rect -1139 -159 -1137 -151
rect -1135 -159 -1133 -151
rect -1070 -159 -1068 -151
rect -1066 -159 -1064 -151
rect -1042 -159 -1040 -151
rect -1038 -159 -1036 -151
rect -984 -159 -982 -151
rect -980 -159 -978 -151
rect -956 -159 -954 -151
rect -952 -159 -950 -151
rect -910 -159 -908 -151
rect -906 -159 -904 -151
rect -882 -159 -880 -151
rect -878 -159 -876 -151
rect -756 -159 -754 -151
rect -752 -159 -750 -151
rect -728 -159 -726 -151
rect -724 -159 -722 -151
rect -660 -159 -658 -151
rect -656 -159 -654 -151
rect -632 -159 -630 -151
rect -628 -159 -626 -151
rect -578 -159 -576 -151
rect -574 -159 -572 -151
rect -550 -159 -548 -151
rect -546 -159 -544 -151
rect -496 -159 -494 -151
rect -492 -159 -490 -151
rect -468 -159 -466 -151
rect -464 -159 -462 -151
rect -1164 -239 -1161 -231
rect -1159 -239 -1156 -231
rect -753 -235 -750 -227
rect -748 -235 -745 -227
rect -1234 -352 -1231 -344
rect -1229 -352 -1226 -344
rect -1167 -350 -1165 -342
rect -1163 -350 -1161 -342
rect -1139 -350 -1137 -342
rect -1135 -350 -1133 -342
rect -1070 -350 -1068 -342
rect -1066 -350 -1064 -342
rect -1042 -350 -1040 -342
rect -1038 -350 -1036 -342
rect -984 -350 -982 -342
rect -980 -350 -978 -342
rect -956 -350 -954 -342
rect -952 -350 -950 -342
rect -910 -350 -908 -342
rect -906 -350 -904 -342
rect -882 -350 -880 -342
rect -878 -350 -876 -342
rect -756 -350 -754 -342
rect -752 -350 -750 -342
rect -728 -350 -726 -342
rect -724 -350 -722 -342
rect -660 -350 -658 -342
rect -656 -350 -654 -342
rect -632 -350 -630 -342
rect -628 -350 -626 -342
rect -578 -350 -576 -342
rect -574 -350 -572 -342
rect -550 -350 -548 -342
rect -546 -350 -544 -342
rect -496 -350 -494 -342
rect -492 -350 -490 -342
rect -468 -350 -466 -342
rect -464 -350 -462 -342
rect -1164 -430 -1161 -422
rect -1159 -430 -1156 -422
rect -753 -426 -750 -418
rect -748 -426 -745 -418
rect -1235 -538 -1232 -530
rect -1230 -538 -1227 -530
rect -1168 -536 -1166 -528
rect -1164 -536 -1162 -528
rect -1140 -536 -1138 -528
rect -1136 -536 -1134 -528
rect -1071 -536 -1069 -528
rect -1067 -536 -1065 -528
rect -1043 -536 -1041 -528
rect -1039 -536 -1037 -528
rect -985 -536 -983 -528
rect -981 -536 -979 -528
rect -957 -536 -955 -528
rect -953 -536 -951 -528
rect -911 -536 -909 -528
rect -907 -536 -905 -528
rect -883 -536 -881 -528
rect -879 -536 -877 -528
rect -757 -536 -755 -528
rect -753 -536 -751 -528
rect -729 -536 -727 -528
rect -725 -536 -723 -528
rect -661 -536 -659 -528
rect -657 -536 -655 -528
rect -633 -536 -631 -528
rect -629 -536 -627 -528
rect -579 -536 -577 -528
rect -575 -536 -573 -528
rect -551 -536 -549 -528
rect -547 -536 -545 -528
rect -497 -536 -495 -528
rect -493 -536 -491 -528
rect -469 -536 -467 -528
rect -465 -536 -463 -528
rect -1165 -616 -1162 -608
rect -1160 -616 -1157 -608
rect -754 -612 -751 -604
rect -749 -612 -746 -604
rect -1218 -709 -1216 -701
rect -1214 -709 -1212 -701
rect -1190 -709 -1188 -701
rect -1186 -709 -1184 -701
rect -1135 -709 -1133 -701
rect -1131 -709 -1129 -701
rect -1107 -709 -1105 -701
rect -1103 -709 -1101 -701
rect -1028 -709 -1026 -701
rect -1024 -709 -1022 -701
rect -1000 -709 -998 -701
rect -996 -709 -994 -701
rect -945 -709 -943 -701
rect -941 -709 -939 -701
rect -917 -709 -915 -701
rect -913 -709 -911 -701
<< metal1 >>
rect -1346 59 -478 63
rect -1346 -129 -1342 59
rect -1286 47 -1282 59
rect -1223 48 -1219 59
rect -1153 49 -1149 59
rect -1056 49 -1052 59
rect -970 49 -966 59
rect -896 49 -892 59
rect -1234 44 -1223 48
rect -1167 45 -1163 49
rect -1159 45 -1153 49
rect -1149 45 -1143 49
rect -1139 45 -1133 49
rect -1238 39 -1234 44
rect -1171 41 -1167 45
rect -1133 41 -1129 45
rect -1157 33 -1143 41
rect -1070 45 -1066 49
rect -1062 45 -1056 49
rect -1052 45 -1046 49
rect -1042 45 -1036 49
rect -1074 41 -1070 45
rect -1036 41 -1032 45
rect -1060 33 -1046 41
rect -984 45 -980 49
rect -976 45 -970 49
rect -966 45 -960 49
rect -956 45 -950 49
rect -988 41 -984 45
rect -950 41 -946 45
rect -974 33 -960 41
rect -910 45 -906 49
rect -902 45 -896 49
rect -892 45 -886 49
rect -882 45 -876 49
rect -914 41 -910 45
rect -876 41 -872 45
rect -819 47 -815 59
rect -742 49 -738 59
rect -646 49 -642 59
rect -564 49 -560 59
rect -482 49 -478 59
rect -756 45 -752 49
rect -748 45 -742 49
rect -738 45 -732 49
rect -728 45 -722 49
rect -900 33 -886 41
rect -1226 21 -1222 31
rect -1187 21 -1169 25
rect -1252 17 -1238 21
rect -1226 17 -1207 21
rect -1226 10 -1222 17
rect -1238 1 -1234 6
rect -1187 3 -1183 21
rect -1153 18 -1149 33
rect -1111 25 -1107 29
rect -1131 21 -1107 25
rect -1086 21 -1072 25
rect -1056 18 -1052 33
rect -1014 25 -1010 29
rect -1034 21 -1010 25
rect -1004 21 -986 25
rect -1004 18 -1000 21
rect -970 18 -966 33
rect -936 25 -932 29
rect -948 21 -932 25
rect -924 21 -912 25
rect -924 18 -920 21
rect -896 18 -892 33
rect -874 21 -864 25
rect -1172 14 -1104 18
rect -1075 14 -1000 18
rect -989 14 -920 18
rect -915 14 -864 18
rect -1172 11 -1168 14
rect -1075 11 -1071 14
rect -989 11 -985 14
rect -915 11 -911 14
rect -868 11 -864 14
rect -855 12 -851 38
rect -760 41 -756 45
rect -722 41 -718 45
rect -746 33 -732 41
rect -660 45 -656 49
rect -652 45 -646 49
rect -642 45 -636 49
rect -632 45 -626 49
rect -664 41 -660 45
rect -626 41 -622 45
rect -650 33 -636 41
rect -578 45 -574 49
rect -570 45 -564 49
rect -560 45 -554 49
rect -550 45 -544 49
rect -582 41 -578 45
rect -544 41 -540 45
rect -568 33 -554 41
rect -496 45 -492 49
rect -488 45 -482 49
rect -478 45 -472 49
rect -468 45 -462 49
rect -500 41 -496 45
rect -462 41 -458 45
rect -486 33 -472 41
rect -776 21 -758 25
rect -776 12 -772 21
rect -742 18 -738 33
rect -700 25 -696 29
rect -720 21 -696 25
rect -676 22 -662 26
rect -646 19 -642 33
rect -604 26 -600 29
rect -624 22 -600 26
rect -592 21 -580 25
rect -592 19 -588 21
rect -855 11 -772 12
rect -1156 7 -1144 11
rect -1059 7 -1047 11
rect -973 7 -961 11
rect -899 7 -887 11
rect -868 8 -772 11
rect -1132 2 -1128 7
rect -1238 -5 -1234 -3
rect -1132 -5 -1128 -2
rect -1035 1 -1031 7
rect -1035 -5 -1031 -3
rect -949 2 -945 7
rect -949 -5 -945 -2
rect -875 1 -871 7
rect -776 3 -772 8
rect -761 14 -692 18
rect -665 15 -588 19
rect -564 18 -560 33
rect -522 25 -518 29
rect -542 21 -518 25
rect -511 21 -498 25
rect -511 18 -507 21
rect -482 18 -478 33
rect -460 21 -450 25
rect -761 11 -757 14
rect -665 12 -661 15
rect -583 14 -507 18
rect -501 14 -450 18
rect -745 7 -733 11
rect -649 8 -637 12
rect -721 1 -717 7
rect -875 -5 -871 -3
rect -721 -5 -717 -3
rect -625 2 -621 8
rect -583 11 -579 14
rect -501 11 -497 14
rect -454 12 -450 14
rect -441 12 -437 38
rect -567 7 -555 11
rect -485 7 -473 11
rect -454 8 -342 12
rect -625 -5 -621 -2
rect -543 2 -539 7
rect -543 -5 -539 -2
rect -461 2 -457 7
rect -461 -5 -457 -2
rect -1331 -9 -457 -5
rect -1301 -19 -1273 -15
rect -1301 -101 -1297 -19
rect -1220 -83 -1216 -9
rect -1134 -16 -1090 -12
rect -1199 -57 -1195 -26
rect -1182 -34 -1168 -30
rect -1164 -34 -1153 -30
rect -1168 -39 -1164 -34
rect -1156 -57 -1152 -47
rect -1134 -57 -1130 -16
rect -1199 -61 -1168 -57
rect -1156 -61 -1130 -57
rect -1156 -68 -1152 -61
rect -1168 -77 -1164 -72
rect -1168 -83 -1164 -81
rect -809 -79 -805 -9
rect -717 -16 -680 -12
rect -788 -53 -784 -20
rect -771 -30 -757 -26
rect -753 -30 -742 -26
rect -757 -35 -753 -30
rect -745 -53 -741 -43
rect -717 -53 -713 -16
rect -788 -57 -757 -53
rect -745 -57 -713 -53
rect -745 -64 -741 -57
rect -757 -73 -753 -68
rect -757 -79 -753 -77
rect -809 -83 -753 -79
rect -1220 -87 -1164 -83
rect -1301 -105 -409 -101
rect -1346 -133 -478 -129
rect -1346 -320 -1342 -133
rect -1286 -145 -1282 -133
rect -1223 -144 -1219 -133
rect -1153 -143 -1149 -133
rect -1056 -143 -1052 -133
rect -970 -143 -966 -133
rect -896 -143 -892 -133
rect -1234 -148 -1223 -144
rect -1167 -147 -1163 -143
rect -1159 -147 -1153 -143
rect -1149 -147 -1143 -143
rect -1139 -147 -1133 -143
rect -1238 -153 -1234 -148
rect -1171 -151 -1167 -147
rect -1133 -151 -1129 -147
rect -1157 -159 -1143 -151
rect -1070 -147 -1066 -143
rect -1062 -147 -1056 -143
rect -1052 -147 -1046 -143
rect -1042 -147 -1036 -143
rect -1074 -151 -1070 -147
rect -1036 -151 -1032 -147
rect -1060 -159 -1046 -151
rect -984 -147 -980 -143
rect -976 -147 -970 -143
rect -966 -147 -960 -143
rect -956 -147 -950 -143
rect -988 -151 -984 -147
rect -950 -151 -946 -147
rect -974 -159 -960 -151
rect -910 -147 -906 -143
rect -902 -147 -896 -143
rect -892 -147 -886 -143
rect -882 -147 -876 -143
rect -914 -151 -910 -147
rect -876 -151 -872 -147
rect -819 -145 -815 -133
rect -742 -143 -738 -133
rect -646 -143 -642 -133
rect -564 -143 -560 -133
rect -482 -143 -478 -133
rect -756 -147 -752 -143
rect -748 -147 -742 -143
rect -738 -147 -732 -143
rect -728 -147 -722 -143
rect -900 -159 -886 -151
rect -1226 -171 -1222 -161
rect -1187 -171 -1169 -167
rect -1252 -175 -1238 -171
rect -1226 -175 -1207 -171
rect -1226 -182 -1222 -175
rect -1238 -191 -1234 -186
rect -1187 -189 -1183 -171
rect -1153 -174 -1149 -159
rect -1111 -167 -1107 -163
rect -1131 -171 -1107 -167
rect -1086 -171 -1072 -167
rect -1056 -174 -1052 -159
rect -1014 -167 -1010 -163
rect -1034 -171 -1010 -167
rect -1004 -171 -986 -167
rect -1004 -174 -1000 -171
rect -970 -174 -966 -159
rect -936 -167 -932 -163
rect -948 -171 -932 -167
rect -924 -171 -912 -167
rect -924 -174 -920 -171
rect -896 -174 -892 -159
rect -874 -171 -864 -167
rect -1172 -178 -1104 -174
rect -1075 -178 -1000 -174
rect -989 -178 -920 -174
rect -915 -178 -864 -174
rect -1172 -181 -1168 -178
rect -1075 -181 -1071 -178
rect -989 -181 -985 -178
rect -915 -181 -911 -178
rect -868 -181 -864 -178
rect -855 -180 -851 -154
rect -760 -151 -756 -147
rect -722 -151 -718 -147
rect -746 -159 -732 -151
rect -660 -147 -656 -143
rect -652 -147 -646 -143
rect -642 -147 -636 -143
rect -632 -147 -626 -143
rect -664 -151 -660 -147
rect -626 -151 -622 -147
rect -650 -159 -636 -151
rect -578 -147 -574 -143
rect -570 -147 -564 -143
rect -560 -147 -554 -143
rect -550 -147 -544 -143
rect -582 -151 -578 -147
rect -544 -151 -540 -147
rect -568 -159 -554 -151
rect -496 -147 -492 -143
rect -488 -147 -482 -143
rect -478 -147 -472 -143
rect -468 -147 -462 -143
rect -500 -151 -496 -147
rect -462 -151 -458 -147
rect -486 -159 -472 -151
rect -776 -171 -758 -167
rect -776 -180 -772 -171
rect -742 -174 -738 -159
rect -700 -167 -696 -163
rect -720 -171 -696 -167
rect -676 -170 -662 -166
rect -646 -173 -642 -159
rect -604 -166 -600 -163
rect -624 -170 -600 -166
rect -592 -171 -580 -167
rect -592 -173 -588 -171
rect -855 -181 -772 -180
rect -1156 -185 -1144 -181
rect -1059 -185 -1047 -181
rect -973 -185 -961 -181
rect -899 -185 -887 -181
rect -868 -184 -772 -181
rect -1132 -190 -1128 -185
rect -1238 -197 -1234 -195
rect -1132 -197 -1128 -194
rect -1035 -191 -1031 -185
rect -1035 -197 -1031 -195
rect -949 -190 -945 -185
rect -949 -197 -945 -194
rect -875 -191 -871 -185
rect -776 -189 -772 -184
rect -761 -178 -692 -174
rect -665 -177 -588 -173
rect -564 -174 -560 -159
rect -522 -167 -518 -163
rect -542 -171 -518 -167
rect -511 -171 -498 -167
rect -511 -174 -507 -171
rect -482 -174 -478 -159
rect -460 -171 -450 -167
rect -761 -181 -757 -178
rect -665 -180 -661 -177
rect -583 -178 -507 -174
rect -501 -178 -450 -174
rect -745 -185 -733 -181
rect -649 -184 -637 -180
rect -721 -191 -717 -185
rect -875 -197 -871 -195
rect -721 -197 -717 -195
rect -625 -190 -621 -184
rect -583 -181 -579 -178
rect -501 -181 -497 -178
rect -454 -180 -450 -178
rect -441 -180 -437 -154
rect -413 -180 -409 -105
rect -567 -185 -555 -181
rect -485 -185 -473 -181
rect -454 -184 -385 -180
rect -625 -197 -621 -194
rect -543 -190 -539 -185
rect -543 -197 -539 -194
rect -461 -190 -457 -185
rect -461 -197 -457 -194
rect -1331 -201 -457 -197
rect -1301 -211 -1273 -207
rect -1301 -289 -1297 -211
rect -1220 -275 -1216 -201
rect -1134 -208 -1090 -204
rect -1199 -249 -1195 -218
rect -1182 -226 -1168 -222
rect -1164 -226 -1153 -222
rect -1168 -231 -1164 -226
rect -1156 -249 -1152 -239
rect -1134 -249 -1130 -208
rect -1199 -253 -1168 -249
rect -1156 -253 -1130 -249
rect -1156 -260 -1152 -253
rect -1168 -269 -1164 -264
rect -1168 -275 -1164 -273
rect -809 -271 -805 -201
rect -717 -208 -680 -204
rect -788 -245 -784 -212
rect -771 -222 -757 -218
rect -753 -222 -742 -218
rect -757 -227 -753 -222
rect -745 -245 -741 -235
rect -717 -245 -713 -208
rect -788 -249 -757 -245
rect -745 -249 -713 -245
rect -745 -256 -741 -249
rect -757 -265 -753 -260
rect -757 -271 -753 -269
rect -809 -275 -753 -271
rect -1220 -279 -1164 -275
rect -1301 -293 -409 -289
rect -1346 -324 -478 -320
rect -1346 -506 -1342 -324
rect -1286 -336 -1282 -324
rect -1223 -335 -1219 -324
rect -1153 -334 -1149 -324
rect -1056 -334 -1052 -324
rect -970 -334 -966 -324
rect -896 -334 -892 -324
rect -1234 -339 -1223 -335
rect -1167 -338 -1163 -334
rect -1159 -338 -1153 -334
rect -1149 -338 -1143 -334
rect -1139 -338 -1133 -334
rect -1238 -344 -1234 -339
rect -1171 -342 -1167 -338
rect -1133 -342 -1129 -338
rect -1157 -350 -1143 -342
rect -1070 -338 -1066 -334
rect -1062 -338 -1056 -334
rect -1052 -338 -1046 -334
rect -1042 -338 -1036 -334
rect -1074 -342 -1070 -338
rect -1036 -342 -1032 -338
rect -1060 -350 -1046 -342
rect -984 -338 -980 -334
rect -976 -338 -970 -334
rect -966 -338 -960 -334
rect -956 -338 -950 -334
rect -988 -342 -984 -338
rect -950 -342 -946 -338
rect -974 -350 -960 -342
rect -910 -338 -906 -334
rect -902 -338 -896 -334
rect -892 -338 -886 -334
rect -882 -338 -876 -334
rect -914 -342 -910 -338
rect -876 -342 -872 -338
rect -819 -336 -815 -324
rect -742 -334 -738 -324
rect -646 -334 -642 -324
rect -564 -334 -560 -324
rect -482 -334 -478 -324
rect -756 -338 -752 -334
rect -748 -338 -742 -334
rect -738 -338 -732 -334
rect -728 -338 -722 -334
rect -900 -350 -886 -342
rect -1226 -362 -1222 -352
rect -1187 -362 -1169 -358
rect -1252 -366 -1238 -362
rect -1226 -366 -1207 -362
rect -1226 -373 -1222 -366
rect -1238 -382 -1234 -377
rect -1187 -380 -1183 -362
rect -1153 -365 -1149 -350
rect -1111 -358 -1107 -354
rect -1131 -362 -1107 -358
rect -1086 -362 -1072 -358
rect -1056 -365 -1052 -350
rect -1014 -358 -1010 -354
rect -1034 -362 -1010 -358
rect -1004 -362 -986 -358
rect -1004 -365 -1000 -362
rect -970 -365 -966 -350
rect -936 -358 -932 -354
rect -948 -362 -932 -358
rect -924 -362 -912 -358
rect -924 -365 -920 -362
rect -896 -365 -892 -350
rect -874 -362 -864 -358
rect -1172 -369 -1104 -365
rect -1075 -369 -1000 -365
rect -989 -369 -920 -365
rect -915 -369 -864 -365
rect -1172 -372 -1168 -369
rect -1075 -372 -1071 -369
rect -989 -372 -985 -369
rect -915 -372 -911 -369
rect -868 -372 -864 -369
rect -855 -371 -851 -345
rect -760 -342 -756 -338
rect -722 -342 -718 -338
rect -746 -350 -732 -342
rect -660 -338 -656 -334
rect -652 -338 -646 -334
rect -642 -338 -636 -334
rect -632 -338 -626 -334
rect -664 -342 -660 -338
rect -626 -342 -622 -338
rect -650 -350 -636 -342
rect -578 -338 -574 -334
rect -570 -338 -564 -334
rect -560 -338 -554 -334
rect -550 -338 -544 -334
rect -582 -342 -578 -338
rect -544 -342 -540 -338
rect -568 -350 -554 -342
rect -496 -338 -492 -334
rect -488 -338 -482 -334
rect -478 -338 -472 -334
rect -468 -338 -462 -334
rect -500 -342 -496 -338
rect -462 -342 -458 -338
rect -486 -350 -472 -342
rect -776 -362 -758 -358
rect -776 -371 -772 -362
rect -742 -365 -738 -350
rect -700 -358 -696 -354
rect -720 -362 -696 -358
rect -676 -361 -662 -357
rect -646 -364 -642 -350
rect -604 -357 -600 -354
rect -624 -361 -600 -357
rect -592 -362 -580 -358
rect -592 -364 -588 -362
rect -855 -372 -772 -371
rect -1156 -376 -1144 -372
rect -1059 -376 -1047 -372
rect -973 -376 -961 -372
rect -899 -376 -887 -372
rect -868 -375 -772 -372
rect -1132 -381 -1128 -376
rect -1238 -388 -1234 -386
rect -1132 -388 -1128 -385
rect -1035 -382 -1031 -376
rect -1035 -388 -1031 -386
rect -949 -381 -945 -376
rect -949 -388 -945 -385
rect -875 -382 -871 -376
rect -776 -380 -772 -375
rect -761 -369 -692 -365
rect -665 -368 -588 -364
rect -564 -365 -560 -350
rect -522 -358 -518 -354
rect -542 -362 -518 -358
rect -511 -362 -498 -358
rect -511 -365 -507 -362
rect -482 -365 -478 -350
rect -460 -362 -450 -358
rect -761 -372 -757 -369
rect -665 -371 -661 -368
rect -583 -369 -507 -365
rect -501 -369 -450 -365
rect -745 -376 -733 -372
rect -649 -375 -637 -371
rect -721 -382 -717 -376
rect -875 -388 -871 -386
rect -721 -388 -717 -386
rect -625 -381 -621 -375
rect -583 -372 -579 -369
rect -501 -372 -497 -369
rect -454 -371 -450 -369
rect -441 -371 -437 -345
rect -413 -371 -409 -293
rect -567 -376 -555 -372
rect -485 -376 -473 -372
rect -454 -375 -385 -371
rect -625 -388 -621 -385
rect -543 -381 -539 -376
rect -543 -388 -539 -385
rect -461 -381 -457 -376
rect -461 -388 -457 -385
rect -1331 -392 -457 -388
rect -1301 -402 -1273 -398
rect -1301 -477 -1297 -402
rect -1220 -466 -1216 -392
rect -1134 -399 -1090 -395
rect -1199 -440 -1195 -409
rect -1182 -417 -1168 -413
rect -1164 -417 -1153 -413
rect -1168 -422 -1164 -417
rect -1156 -440 -1152 -430
rect -1134 -440 -1130 -399
rect -1199 -444 -1168 -440
rect -1156 -444 -1130 -440
rect -1156 -451 -1152 -444
rect -1168 -460 -1164 -455
rect -1168 -466 -1164 -464
rect -809 -462 -805 -392
rect -717 -399 -680 -395
rect -788 -436 -784 -403
rect -771 -413 -757 -409
rect -753 -413 -742 -409
rect -757 -418 -753 -413
rect -745 -436 -741 -426
rect -717 -436 -713 -399
rect -788 -440 -757 -436
rect -745 -440 -713 -436
rect -745 -447 -741 -440
rect -757 -456 -753 -451
rect -757 -462 -753 -460
rect -809 -466 -753 -462
rect -1220 -470 -1164 -466
rect -1301 -481 -388 -477
rect -1356 -510 -479 -506
rect -1346 -675 -1342 -510
rect -1287 -522 -1283 -510
rect -1224 -521 -1220 -510
rect -1154 -520 -1150 -510
rect -1057 -520 -1053 -510
rect -971 -520 -967 -510
rect -897 -520 -893 -510
rect -1235 -525 -1224 -521
rect -1168 -524 -1164 -520
rect -1160 -524 -1154 -520
rect -1150 -524 -1144 -520
rect -1140 -524 -1134 -520
rect -1239 -530 -1235 -525
rect -1172 -528 -1168 -524
rect -1134 -528 -1130 -524
rect -1158 -536 -1144 -528
rect -1071 -524 -1067 -520
rect -1063 -524 -1057 -520
rect -1053 -524 -1047 -520
rect -1043 -524 -1037 -520
rect -1075 -528 -1071 -524
rect -1037 -528 -1033 -524
rect -1061 -536 -1047 -528
rect -985 -524 -981 -520
rect -977 -524 -971 -520
rect -967 -524 -961 -520
rect -957 -524 -951 -520
rect -989 -528 -985 -524
rect -951 -528 -947 -524
rect -975 -536 -961 -528
rect -911 -524 -907 -520
rect -903 -524 -897 -520
rect -893 -524 -887 -520
rect -883 -524 -877 -520
rect -915 -528 -911 -524
rect -877 -528 -873 -524
rect -820 -522 -816 -510
rect -743 -520 -739 -510
rect -647 -520 -643 -510
rect -565 -520 -561 -510
rect -483 -520 -479 -510
rect -757 -524 -753 -520
rect -749 -524 -743 -520
rect -739 -524 -733 -520
rect -729 -524 -723 -520
rect -901 -536 -887 -528
rect -1227 -548 -1223 -538
rect -1188 -548 -1170 -544
rect -1253 -552 -1239 -548
rect -1227 -552 -1208 -548
rect -1227 -559 -1223 -552
rect -1239 -568 -1235 -563
rect -1188 -566 -1184 -548
rect -1154 -551 -1150 -536
rect -1112 -544 -1108 -540
rect -1132 -548 -1108 -544
rect -1087 -548 -1073 -544
rect -1057 -551 -1053 -536
rect -1015 -544 -1011 -540
rect -1035 -548 -1011 -544
rect -1005 -548 -987 -544
rect -1005 -551 -1001 -548
rect -971 -551 -967 -536
rect -937 -544 -933 -540
rect -949 -548 -933 -544
rect -925 -548 -913 -544
rect -925 -551 -921 -548
rect -897 -551 -893 -536
rect -875 -548 -865 -544
rect -1173 -555 -1105 -551
rect -1076 -555 -1001 -551
rect -990 -555 -921 -551
rect -916 -555 -865 -551
rect -1173 -558 -1169 -555
rect -1076 -558 -1072 -555
rect -990 -558 -986 -555
rect -916 -558 -912 -555
rect -869 -558 -865 -555
rect -856 -557 -852 -531
rect -761 -528 -757 -524
rect -723 -528 -719 -524
rect -747 -536 -733 -528
rect -661 -524 -657 -520
rect -653 -524 -647 -520
rect -643 -524 -637 -520
rect -633 -524 -627 -520
rect -665 -528 -661 -524
rect -627 -528 -623 -524
rect -651 -536 -637 -528
rect -579 -524 -575 -520
rect -571 -524 -565 -520
rect -561 -524 -555 -520
rect -551 -524 -545 -520
rect -583 -528 -579 -524
rect -545 -528 -541 -524
rect -569 -536 -555 -528
rect -497 -524 -493 -520
rect -489 -524 -483 -520
rect -479 -524 -473 -520
rect -469 -524 -463 -520
rect -501 -528 -497 -524
rect -463 -528 -459 -524
rect -487 -536 -473 -528
rect -777 -548 -759 -544
rect -777 -557 -773 -548
rect -743 -551 -739 -536
rect -701 -544 -697 -540
rect -721 -548 -697 -544
rect -677 -547 -663 -543
rect -647 -550 -643 -536
rect -605 -543 -601 -540
rect -625 -547 -601 -543
rect -593 -548 -581 -544
rect -593 -550 -589 -548
rect -856 -558 -773 -557
rect -1157 -562 -1145 -558
rect -1060 -562 -1048 -558
rect -974 -562 -962 -558
rect -900 -562 -888 -558
rect -869 -561 -773 -558
rect -1133 -567 -1129 -562
rect -1239 -574 -1235 -572
rect -1133 -574 -1129 -571
rect -1036 -568 -1032 -562
rect -1036 -574 -1032 -572
rect -950 -567 -946 -562
rect -950 -574 -946 -571
rect -876 -568 -872 -562
rect -777 -566 -773 -561
rect -762 -555 -693 -551
rect -666 -554 -589 -550
rect -565 -551 -561 -536
rect -523 -544 -519 -540
rect -543 -548 -519 -544
rect -512 -548 -499 -544
rect -512 -551 -508 -548
rect -483 -551 -479 -536
rect -461 -548 -451 -544
rect -762 -558 -758 -555
rect -666 -557 -662 -554
rect -584 -555 -508 -551
rect -502 -555 -451 -551
rect -746 -562 -734 -558
rect -650 -561 -638 -557
rect -722 -568 -718 -562
rect -876 -574 -872 -572
rect -722 -574 -718 -572
rect -626 -567 -622 -561
rect -584 -558 -580 -555
rect -502 -558 -498 -555
rect -455 -557 -451 -555
rect -442 -557 -438 -531
rect -392 -557 -388 -481
rect -568 -562 -556 -558
rect -486 -562 -474 -558
rect -455 -561 -384 -557
rect -626 -574 -622 -571
rect -544 -567 -540 -562
rect -544 -574 -540 -571
rect -462 -567 -458 -562
rect -462 -574 -458 -571
rect -1331 -578 -458 -574
rect -1297 -588 -1274 -584
rect -1297 -648 -1293 -588
rect -1221 -652 -1217 -578
rect -1135 -585 -1091 -581
rect -1200 -626 -1196 -595
rect -1183 -603 -1169 -599
rect -1165 -603 -1154 -599
rect -1169 -608 -1165 -603
rect -1157 -626 -1153 -616
rect -1135 -626 -1131 -585
rect -1200 -630 -1169 -626
rect -1157 -630 -1131 -626
rect -1157 -637 -1153 -630
rect -1169 -646 -1165 -641
rect -1169 -652 -1165 -650
rect -810 -648 -806 -578
rect -718 -585 -681 -581
rect -789 -622 -785 -589
rect -772 -599 -758 -595
rect -754 -599 -743 -595
rect -758 -604 -754 -599
rect -746 -622 -742 -612
rect -718 -622 -714 -585
rect -789 -626 -758 -622
rect -746 -626 -714 -622
rect -746 -633 -742 -626
rect -758 -642 -754 -637
rect -758 -648 -754 -646
rect -810 -652 -754 -648
rect -1221 -656 -1165 -652
rect -392 -659 -388 -561
rect -1049 -663 -388 -659
rect -1346 -679 -927 -675
rect -1204 -693 -1200 -679
rect -1121 -693 -1117 -679
rect -1014 -693 -1010 -679
rect -931 -693 -927 -679
rect -1218 -697 -1214 -693
rect -1210 -697 -1204 -693
rect -1200 -697 -1194 -693
rect -1190 -697 -1184 -693
rect -1222 -701 -1218 -697
rect -1184 -701 -1180 -697
rect -1208 -709 -1194 -701
rect -1135 -697 -1131 -693
rect -1127 -697 -1121 -693
rect -1117 -697 -1111 -693
rect -1107 -697 -1101 -693
rect -1139 -701 -1135 -697
rect -1101 -701 -1097 -697
rect -1125 -709 -1111 -701
rect -1028 -697 -1024 -693
rect -1020 -697 -1014 -693
rect -1010 -697 -1004 -693
rect -1000 -697 -994 -693
rect -1032 -701 -1028 -697
rect -994 -701 -990 -697
rect -945 -697 -941 -693
rect -937 -697 -931 -693
rect -927 -697 -921 -693
rect -917 -697 -911 -693
rect -1018 -709 -1004 -701
rect -1235 -721 -1220 -717
rect -1204 -724 -1200 -709
rect -1182 -721 -1165 -717
rect -1148 -721 -1137 -717
rect -1293 -728 -1200 -724
rect -1169 -724 -1165 -721
rect -1121 -724 -1117 -709
rect -1099 -721 -1086 -717
rect -1049 -721 -1030 -717
rect -1014 -724 -1010 -709
rect -965 -717 -961 -703
rect -949 -701 -945 -697
rect -911 -701 -907 -697
rect -935 -709 -921 -701
rect -992 -721 -975 -717
rect -965 -721 -947 -717
rect -1169 -728 -1117 -724
rect -1069 -728 -1010 -724
rect -979 -724 -975 -721
rect -931 -724 -927 -709
rect -392 -717 -388 -663
rect -346 -663 -342 8
rect -909 -721 -388 -717
rect -979 -728 -927 -724
rect -1223 -731 -1219 -728
rect -1140 -731 -1136 -728
rect -1033 -731 -1029 -728
rect -1207 -735 -1195 -731
rect -1124 -735 -1112 -731
rect -1017 -735 -1005 -731
rect -1183 -741 -1179 -735
rect -1183 -747 -1179 -745
rect -1100 -741 -1096 -735
rect -1100 -747 -1096 -745
rect -993 -741 -989 -735
rect -959 -737 -955 -728
rect -950 -731 -946 -728
rect -934 -735 -922 -731
rect -910 -741 -906 -735
rect -993 -747 -989 -745
rect -910 -747 -906 -745
rect -1331 -751 -906 -747
<< metal2 >>
rect -1320 66 -600 70
rect -1335 -197 -1331 -9
rect -1335 -388 -1331 -201
rect -1335 -574 -1331 -392
rect -1335 -747 -1331 -578
rect -1320 -122 -1316 66
rect -1286 -30 -1282 43
rect -1256 21 -1252 66
rect -1196 53 -1010 57
rect -1196 21 -1192 53
rect -1111 33 -1107 53
rect -1014 33 -1010 53
rect -936 55 -851 59
rect -936 33 -932 55
rect -855 43 -851 55
rect -1203 17 -1192 21
rect -860 21 -832 25
rect -1199 -1 -1187 3
rect -1199 -15 -1195 -1
rect -1269 -19 -1195 -15
rect -1199 -22 -1195 -19
rect -1104 -25 -1100 14
rect -1090 -12 -1086 21
rect -836 -25 -832 21
rect -1104 -29 -832 -25
rect -819 -26 -815 43
rect -700 33 -696 66
rect -604 33 -600 66
rect -522 54 -437 58
rect -522 33 -518 54
rect -441 42 -437 54
rect -788 -1 -776 3
rect -788 -16 -784 -1
rect -692 -23 -688 14
rect -680 -12 -676 22
rect -446 21 -424 25
rect -428 -23 -424 21
rect -819 -30 -775 -26
rect -692 -27 -424 -23
rect -1286 -34 -1186 -30
rect -1320 -126 -600 -122
rect -1320 -313 -1316 -126
rect -1286 -222 -1282 -149
rect -1256 -171 -1252 -126
rect -1196 -139 -1010 -135
rect -1196 -171 -1192 -139
rect -1111 -159 -1107 -139
rect -1014 -159 -1010 -139
rect -936 -137 -851 -133
rect -936 -159 -932 -137
rect -855 -149 -851 -137
rect -1203 -175 -1192 -171
rect -860 -171 -832 -167
rect -1199 -193 -1187 -189
rect -1199 -207 -1195 -193
rect -1269 -211 -1195 -207
rect -1199 -214 -1195 -211
rect -1104 -217 -1100 -178
rect -1090 -204 -1086 -171
rect -836 -217 -832 -171
rect -1104 -221 -832 -217
rect -819 -218 -815 -149
rect -700 -159 -696 -126
rect -604 -159 -600 -126
rect -522 -138 -437 -134
rect -522 -159 -518 -138
rect -441 -150 -437 -138
rect -788 -193 -776 -189
rect -788 -208 -784 -193
rect -692 -215 -688 -178
rect -680 -204 -676 -170
rect -446 -171 -424 -167
rect -428 -215 -424 -171
rect -819 -222 -775 -218
rect -692 -219 -424 -215
rect -1286 -226 -1186 -222
rect -1320 -317 -600 -313
rect -1320 -499 -1316 -317
rect -1286 -413 -1282 -340
rect -1256 -362 -1252 -317
rect -1196 -330 -1010 -326
rect -1196 -362 -1192 -330
rect -1111 -350 -1107 -330
rect -1014 -350 -1010 -330
rect -936 -328 -851 -324
rect -936 -350 -932 -328
rect -855 -340 -851 -328
rect -1203 -366 -1192 -362
rect -860 -362 -832 -358
rect -1199 -384 -1187 -380
rect -1199 -398 -1195 -384
rect -1269 -402 -1195 -398
rect -1199 -405 -1195 -402
rect -1104 -408 -1100 -369
rect -1090 -395 -1086 -362
rect -836 -408 -832 -362
rect -1104 -412 -832 -408
rect -819 -409 -815 -340
rect -700 -350 -696 -317
rect -604 -350 -600 -317
rect -522 -329 -437 -325
rect -522 -350 -518 -329
rect -441 -341 -437 -329
rect -788 -384 -776 -380
rect -788 -399 -784 -384
rect -692 -406 -688 -369
rect -680 -395 -676 -361
rect -446 -362 -424 -358
rect -428 -406 -424 -362
rect -819 -413 -775 -409
rect -692 -410 -424 -406
rect -1286 -417 -1186 -413
rect -1320 -503 -601 -499
rect -1320 -607 -1316 -503
rect -1287 -599 -1283 -526
rect -1257 -548 -1253 -503
rect -1197 -516 -1011 -512
rect -1197 -548 -1193 -516
rect -1112 -536 -1108 -516
rect -1015 -536 -1011 -516
rect -937 -514 -852 -510
rect -937 -536 -933 -514
rect -856 -526 -852 -514
rect -1204 -552 -1193 -548
rect -861 -548 -833 -544
rect -1200 -570 -1188 -566
rect -1200 -584 -1196 -570
rect -1269 -588 -1196 -584
rect -1200 -591 -1196 -588
rect -1105 -594 -1101 -555
rect -1091 -581 -1087 -548
rect -837 -594 -833 -548
rect -1105 -598 -833 -594
rect -820 -595 -816 -526
rect -701 -536 -697 -503
rect -605 -536 -601 -503
rect -523 -515 -438 -511
rect -523 -536 -519 -515
rect -442 -527 -438 -515
rect -789 -570 -777 -566
rect -789 -585 -785 -570
rect -693 -592 -689 -555
rect -681 -581 -677 -547
rect -447 -548 -425 -544
rect -429 -592 -425 -548
rect -820 -599 -776 -595
rect -693 -596 -425 -592
rect -1287 -603 -1187 -599
rect -1297 -724 -1293 -652
rect -1239 -672 -1069 -668
rect -1239 -717 -1235 -672
rect -1335 -806 -1331 -751
rect -1152 -777 -1148 -721
rect -1086 -756 -1082 -721
rect -1073 -724 -1069 -672
rect -1053 -717 -1049 -663
rect -965 -667 -346 -663
rect -965 -699 -961 -667
rect -959 -756 -955 -741
rect -1086 -760 -955 -756
rect -824 -777 -820 -667
rect -1152 -781 -820 -777
<< ntransistor >>
rect -1231 6 -1229 10
rect -1165 7 -1163 11
rect -1137 7 -1135 11
rect -1068 7 -1066 11
rect -1040 7 -1038 11
rect -982 7 -980 11
rect -954 7 -952 11
rect -908 7 -906 11
rect -880 7 -878 11
rect -754 7 -752 11
rect -726 7 -724 11
rect -658 8 -656 12
rect -630 8 -628 12
rect -576 7 -574 11
rect -548 7 -546 11
rect -494 7 -492 11
rect -466 7 -464 11
rect -750 -68 -748 -64
rect -1161 -72 -1159 -68
rect -1231 -186 -1229 -182
rect -1165 -185 -1163 -181
rect -1137 -185 -1135 -181
rect -1068 -185 -1066 -181
rect -1040 -185 -1038 -181
rect -982 -185 -980 -181
rect -954 -185 -952 -181
rect -908 -185 -906 -181
rect -880 -185 -878 -181
rect -754 -185 -752 -181
rect -726 -185 -724 -181
rect -658 -184 -656 -180
rect -630 -184 -628 -180
rect -576 -185 -574 -181
rect -548 -185 -546 -181
rect -494 -185 -492 -181
rect -466 -185 -464 -181
rect -750 -260 -748 -256
rect -1161 -264 -1159 -260
rect -1231 -377 -1229 -373
rect -1165 -376 -1163 -372
rect -1137 -376 -1135 -372
rect -1068 -376 -1066 -372
rect -1040 -376 -1038 -372
rect -982 -376 -980 -372
rect -954 -376 -952 -372
rect -908 -376 -906 -372
rect -880 -376 -878 -372
rect -754 -376 -752 -372
rect -726 -376 -724 -372
rect -658 -375 -656 -371
rect -630 -375 -628 -371
rect -576 -376 -574 -372
rect -548 -376 -546 -372
rect -494 -376 -492 -372
rect -466 -376 -464 -372
rect -750 -451 -748 -447
rect -1161 -455 -1159 -451
rect -1232 -563 -1230 -559
rect -1166 -562 -1164 -558
rect -1138 -562 -1136 -558
rect -1069 -562 -1067 -558
rect -1041 -562 -1039 -558
rect -983 -562 -981 -558
rect -955 -562 -953 -558
rect -909 -562 -907 -558
rect -881 -562 -879 -558
rect -755 -562 -753 -558
rect -727 -562 -725 -558
rect -659 -561 -657 -557
rect -631 -561 -629 -557
rect -577 -562 -575 -558
rect -549 -562 -547 -558
rect -495 -562 -493 -558
rect -467 -562 -465 -558
rect -751 -637 -749 -633
rect -1162 -641 -1160 -637
rect -1216 -735 -1214 -731
rect -1188 -735 -1186 -731
rect -1133 -735 -1131 -731
rect -1105 -735 -1103 -731
rect -1026 -735 -1024 -731
rect -998 -735 -996 -731
rect -943 -735 -941 -731
rect -915 -735 -913 -731
<< ptransistor >>
rect -1231 31 -1229 39
rect -1165 33 -1163 41
rect -1137 33 -1135 41
rect -1068 33 -1066 41
rect -1040 33 -1038 41
rect -982 33 -980 41
rect -954 33 -952 41
rect -908 33 -906 41
rect -880 33 -878 41
rect -754 33 -752 41
rect -726 33 -724 41
rect -658 33 -656 41
rect -630 33 -628 41
rect -576 33 -574 41
rect -548 33 -546 41
rect -494 33 -492 41
rect -466 33 -464 41
rect -1161 -47 -1159 -39
rect -750 -43 -748 -35
rect -1231 -161 -1229 -153
rect -1165 -159 -1163 -151
rect -1137 -159 -1135 -151
rect -1068 -159 -1066 -151
rect -1040 -159 -1038 -151
rect -982 -159 -980 -151
rect -954 -159 -952 -151
rect -908 -159 -906 -151
rect -880 -159 -878 -151
rect -754 -159 -752 -151
rect -726 -159 -724 -151
rect -658 -159 -656 -151
rect -630 -159 -628 -151
rect -576 -159 -574 -151
rect -548 -159 -546 -151
rect -494 -159 -492 -151
rect -466 -159 -464 -151
rect -1161 -239 -1159 -231
rect -750 -235 -748 -227
rect -1231 -352 -1229 -344
rect -1165 -350 -1163 -342
rect -1137 -350 -1135 -342
rect -1068 -350 -1066 -342
rect -1040 -350 -1038 -342
rect -982 -350 -980 -342
rect -954 -350 -952 -342
rect -908 -350 -906 -342
rect -880 -350 -878 -342
rect -754 -350 -752 -342
rect -726 -350 -724 -342
rect -658 -350 -656 -342
rect -630 -350 -628 -342
rect -576 -350 -574 -342
rect -548 -350 -546 -342
rect -494 -350 -492 -342
rect -466 -350 -464 -342
rect -1161 -430 -1159 -422
rect -750 -426 -748 -418
rect -1232 -538 -1230 -530
rect -1166 -536 -1164 -528
rect -1138 -536 -1136 -528
rect -1069 -536 -1067 -528
rect -1041 -536 -1039 -528
rect -983 -536 -981 -528
rect -955 -536 -953 -528
rect -909 -536 -907 -528
rect -881 -536 -879 -528
rect -755 -536 -753 -528
rect -727 -536 -725 -528
rect -659 -536 -657 -528
rect -631 -536 -629 -528
rect -577 -536 -575 -528
rect -549 -536 -547 -528
rect -495 -536 -493 -528
rect -467 -536 -465 -528
rect -1162 -616 -1160 -608
rect -751 -612 -749 -604
rect -1216 -709 -1214 -701
rect -1188 -709 -1186 -701
rect -1133 -709 -1131 -701
rect -1105 -709 -1103 -701
rect -1026 -709 -1024 -701
rect -998 -709 -996 -701
rect -943 -709 -941 -701
rect -915 -709 -913 -701
<< polycontact >>
rect -1238 17 -1234 21
rect -1169 21 -1165 25
rect -1135 21 -1131 25
rect -1072 21 -1068 25
rect -1038 21 -1034 25
rect -986 21 -982 25
rect -952 21 -948 25
rect -912 21 -908 25
rect -878 21 -874 25
rect -758 21 -754 25
rect -724 21 -720 25
rect -662 22 -658 26
rect -628 22 -624 26
rect -580 21 -576 25
rect -546 21 -542 25
rect -498 21 -494 25
rect -464 21 -460 25
rect -1168 -61 -1164 -57
rect -757 -57 -753 -53
rect -1238 -175 -1234 -171
rect -1169 -171 -1165 -167
rect -1135 -171 -1131 -167
rect -1072 -171 -1068 -167
rect -1038 -171 -1034 -167
rect -986 -171 -982 -167
rect -952 -171 -948 -167
rect -912 -171 -908 -167
rect -878 -171 -874 -167
rect -758 -171 -754 -167
rect -724 -171 -720 -167
rect -662 -170 -658 -166
rect -628 -170 -624 -166
rect -580 -171 -576 -167
rect -546 -171 -542 -167
rect -498 -171 -494 -167
rect -464 -171 -460 -167
rect -1168 -253 -1164 -249
rect -757 -249 -753 -245
rect -1238 -366 -1234 -362
rect -1169 -362 -1165 -358
rect -1135 -362 -1131 -358
rect -1072 -362 -1068 -358
rect -1038 -362 -1034 -358
rect -986 -362 -982 -358
rect -952 -362 -948 -358
rect -912 -362 -908 -358
rect -878 -362 -874 -358
rect -758 -362 -754 -358
rect -724 -362 -720 -358
rect -662 -361 -658 -357
rect -628 -361 -624 -357
rect -580 -362 -576 -358
rect -546 -362 -542 -358
rect -498 -362 -494 -358
rect -464 -362 -460 -358
rect -1168 -444 -1164 -440
rect -757 -440 -753 -436
rect -1239 -552 -1235 -548
rect -1170 -548 -1166 -544
rect -1136 -548 -1132 -544
rect -1073 -548 -1069 -544
rect -1039 -548 -1035 -544
rect -987 -548 -983 -544
rect -953 -548 -949 -544
rect -913 -548 -909 -544
rect -879 -548 -875 -544
rect -759 -548 -755 -544
rect -725 -548 -721 -544
rect -663 -547 -659 -543
rect -629 -547 -625 -543
rect -581 -548 -577 -544
rect -547 -548 -543 -544
rect -499 -548 -495 -544
rect -465 -548 -461 -544
rect -1169 -630 -1165 -626
rect -758 -626 -754 -622
rect -1220 -721 -1216 -717
rect -1186 -721 -1182 -717
rect -1137 -721 -1133 -717
rect -1103 -721 -1099 -717
rect -1030 -721 -1026 -717
rect -996 -721 -992 -717
rect -947 -721 -943 -717
rect -913 -721 -909 -717
<< ndcontact >>
rect -1238 6 -1234 10
rect -1226 6 -1222 10
rect -1172 7 -1168 11
rect -1160 7 -1156 11
rect -1144 7 -1140 11
rect -1132 7 -1128 11
rect -1075 7 -1071 11
rect -1063 7 -1059 11
rect -1047 7 -1043 11
rect -1035 7 -1031 11
rect -989 7 -985 11
rect -977 7 -973 11
rect -961 7 -957 11
rect -949 7 -945 11
rect -915 7 -911 11
rect -903 7 -899 11
rect -887 7 -883 11
rect -875 7 -871 11
rect -761 7 -757 11
rect -749 7 -745 11
rect -733 7 -729 11
rect -721 7 -717 11
rect -665 8 -661 12
rect -653 8 -649 12
rect -637 8 -633 12
rect -625 8 -621 12
rect -583 7 -579 11
rect -571 7 -567 11
rect -555 7 -551 11
rect -543 7 -539 11
rect -501 7 -497 11
rect -489 7 -485 11
rect -473 7 -469 11
rect -461 7 -457 11
rect -757 -68 -753 -64
rect -745 -68 -741 -64
rect -1168 -72 -1164 -68
rect -1156 -72 -1152 -68
rect -1238 -186 -1234 -182
rect -1226 -186 -1222 -182
rect -1172 -185 -1168 -181
rect -1160 -185 -1156 -181
rect -1144 -185 -1140 -181
rect -1132 -185 -1128 -181
rect -1075 -185 -1071 -181
rect -1063 -185 -1059 -181
rect -1047 -185 -1043 -181
rect -1035 -185 -1031 -181
rect -989 -185 -985 -181
rect -977 -185 -973 -181
rect -961 -185 -957 -181
rect -949 -185 -945 -181
rect -915 -185 -911 -181
rect -903 -185 -899 -181
rect -887 -185 -883 -181
rect -875 -185 -871 -181
rect -761 -185 -757 -181
rect -749 -185 -745 -181
rect -733 -185 -729 -181
rect -721 -185 -717 -181
rect -665 -184 -661 -180
rect -653 -184 -649 -180
rect -637 -184 -633 -180
rect -625 -184 -621 -180
rect -583 -185 -579 -181
rect -571 -185 -567 -181
rect -555 -185 -551 -181
rect -543 -185 -539 -181
rect -501 -185 -497 -181
rect -489 -185 -485 -181
rect -473 -185 -469 -181
rect -461 -185 -457 -181
rect -757 -260 -753 -256
rect -745 -260 -741 -256
rect -1168 -264 -1164 -260
rect -1156 -264 -1152 -260
rect -1238 -377 -1234 -373
rect -1226 -377 -1222 -373
rect -1172 -376 -1168 -372
rect -1160 -376 -1156 -372
rect -1144 -376 -1140 -372
rect -1132 -376 -1128 -372
rect -1075 -376 -1071 -372
rect -1063 -376 -1059 -372
rect -1047 -376 -1043 -372
rect -1035 -376 -1031 -372
rect -989 -376 -985 -372
rect -977 -376 -973 -372
rect -961 -376 -957 -372
rect -949 -376 -945 -372
rect -915 -376 -911 -372
rect -903 -376 -899 -372
rect -887 -376 -883 -372
rect -875 -376 -871 -372
rect -761 -376 -757 -372
rect -749 -376 -745 -372
rect -733 -376 -729 -372
rect -721 -376 -717 -372
rect -665 -375 -661 -371
rect -653 -375 -649 -371
rect -637 -375 -633 -371
rect -625 -375 -621 -371
rect -583 -376 -579 -372
rect -571 -376 -567 -372
rect -555 -376 -551 -372
rect -543 -376 -539 -372
rect -501 -376 -497 -372
rect -489 -376 -485 -372
rect -473 -376 -469 -372
rect -461 -376 -457 -372
rect -757 -451 -753 -447
rect -745 -451 -741 -447
rect -1168 -455 -1164 -451
rect -1156 -455 -1152 -451
rect -1239 -563 -1235 -559
rect -1227 -563 -1223 -559
rect -1173 -562 -1169 -558
rect -1161 -562 -1157 -558
rect -1145 -562 -1141 -558
rect -1133 -562 -1129 -558
rect -1076 -562 -1072 -558
rect -1064 -562 -1060 -558
rect -1048 -562 -1044 -558
rect -1036 -562 -1032 -558
rect -990 -562 -986 -558
rect -978 -562 -974 -558
rect -962 -562 -958 -558
rect -950 -562 -946 -558
rect -916 -562 -912 -558
rect -904 -562 -900 -558
rect -888 -562 -884 -558
rect -876 -562 -872 -558
rect -762 -562 -758 -558
rect -750 -562 -746 -558
rect -734 -562 -730 -558
rect -722 -562 -718 -558
rect -666 -561 -662 -557
rect -654 -561 -650 -557
rect -638 -561 -634 -557
rect -626 -561 -622 -557
rect -584 -562 -580 -558
rect -572 -562 -568 -558
rect -556 -562 -552 -558
rect -544 -562 -540 -558
rect -502 -562 -498 -558
rect -490 -562 -486 -558
rect -474 -562 -470 -558
rect -462 -562 -458 -558
rect -758 -637 -754 -633
rect -746 -637 -742 -633
rect -1169 -641 -1165 -637
rect -1157 -641 -1153 -637
rect -1223 -735 -1219 -731
rect -1211 -735 -1207 -731
rect -1195 -735 -1191 -731
rect -1183 -735 -1179 -731
rect -1140 -735 -1136 -731
rect -1128 -735 -1124 -731
rect -1112 -735 -1108 -731
rect -1100 -735 -1096 -731
rect -1033 -735 -1029 -731
rect -1021 -735 -1017 -731
rect -1005 -735 -1001 -731
rect -993 -735 -989 -731
rect -950 -735 -946 -731
rect -938 -735 -934 -731
rect -922 -735 -918 -731
rect -910 -735 -906 -731
<< pdcontact >>
rect -1238 31 -1234 39
rect -1226 31 -1222 39
rect -1171 33 -1167 41
rect -1161 33 -1157 41
rect -1143 33 -1139 41
rect -1133 33 -1129 41
rect -1074 33 -1070 41
rect -1064 33 -1060 41
rect -1046 33 -1042 41
rect -1036 33 -1032 41
rect -988 33 -984 41
rect -978 33 -974 41
rect -960 33 -956 41
rect -950 33 -946 41
rect -914 33 -910 41
rect -904 33 -900 41
rect -886 33 -882 41
rect -876 33 -872 41
rect -760 33 -756 41
rect -750 33 -746 41
rect -732 33 -728 41
rect -722 33 -718 41
rect -664 33 -660 41
rect -654 33 -650 41
rect -636 33 -632 41
rect -626 33 -622 41
rect -582 33 -578 41
rect -572 33 -568 41
rect -554 33 -550 41
rect -544 33 -540 41
rect -500 33 -496 41
rect -490 33 -486 41
rect -472 33 -468 41
rect -462 33 -458 41
rect -1168 -47 -1164 -39
rect -1156 -47 -1152 -39
rect -757 -43 -753 -35
rect -745 -43 -741 -35
rect -1238 -161 -1234 -153
rect -1226 -161 -1222 -153
rect -1171 -159 -1167 -151
rect -1161 -159 -1157 -151
rect -1143 -159 -1139 -151
rect -1133 -159 -1129 -151
rect -1074 -159 -1070 -151
rect -1064 -159 -1060 -151
rect -1046 -159 -1042 -151
rect -1036 -159 -1032 -151
rect -988 -159 -984 -151
rect -978 -159 -974 -151
rect -960 -159 -956 -151
rect -950 -159 -946 -151
rect -914 -159 -910 -151
rect -904 -159 -900 -151
rect -886 -159 -882 -151
rect -876 -159 -872 -151
rect -760 -159 -756 -151
rect -750 -159 -746 -151
rect -732 -159 -728 -151
rect -722 -159 -718 -151
rect -664 -159 -660 -151
rect -654 -159 -650 -151
rect -636 -159 -632 -151
rect -626 -159 -622 -151
rect -582 -159 -578 -151
rect -572 -159 -568 -151
rect -554 -159 -550 -151
rect -544 -159 -540 -151
rect -500 -159 -496 -151
rect -490 -159 -486 -151
rect -472 -159 -468 -151
rect -462 -159 -458 -151
rect -1168 -239 -1164 -231
rect -1156 -239 -1152 -231
rect -757 -235 -753 -227
rect -745 -235 -741 -227
rect -1238 -352 -1234 -344
rect -1226 -352 -1222 -344
rect -1171 -350 -1167 -342
rect -1161 -350 -1157 -342
rect -1143 -350 -1139 -342
rect -1133 -350 -1129 -342
rect -1074 -350 -1070 -342
rect -1064 -350 -1060 -342
rect -1046 -350 -1042 -342
rect -1036 -350 -1032 -342
rect -988 -350 -984 -342
rect -978 -350 -974 -342
rect -960 -350 -956 -342
rect -950 -350 -946 -342
rect -914 -350 -910 -342
rect -904 -350 -900 -342
rect -886 -350 -882 -342
rect -876 -350 -872 -342
rect -760 -350 -756 -342
rect -750 -350 -746 -342
rect -732 -350 -728 -342
rect -722 -350 -718 -342
rect -664 -350 -660 -342
rect -654 -350 -650 -342
rect -636 -350 -632 -342
rect -626 -350 -622 -342
rect -582 -350 -578 -342
rect -572 -350 -568 -342
rect -554 -350 -550 -342
rect -544 -350 -540 -342
rect -500 -350 -496 -342
rect -490 -350 -486 -342
rect -472 -350 -468 -342
rect -462 -350 -458 -342
rect -1168 -430 -1164 -422
rect -1156 -430 -1152 -422
rect -757 -426 -753 -418
rect -745 -426 -741 -418
rect -1239 -538 -1235 -530
rect -1227 -538 -1223 -530
rect -1172 -536 -1168 -528
rect -1162 -536 -1158 -528
rect -1144 -536 -1140 -528
rect -1134 -536 -1130 -528
rect -1075 -536 -1071 -528
rect -1065 -536 -1061 -528
rect -1047 -536 -1043 -528
rect -1037 -536 -1033 -528
rect -989 -536 -985 -528
rect -979 -536 -975 -528
rect -961 -536 -957 -528
rect -951 -536 -947 -528
rect -915 -536 -911 -528
rect -905 -536 -901 -528
rect -887 -536 -883 -528
rect -877 -536 -873 -528
rect -761 -536 -757 -528
rect -751 -536 -747 -528
rect -733 -536 -729 -528
rect -723 -536 -719 -528
rect -665 -536 -661 -528
rect -655 -536 -651 -528
rect -637 -536 -633 -528
rect -627 -536 -623 -528
rect -583 -536 -579 -528
rect -573 -536 -569 -528
rect -555 -536 -551 -528
rect -545 -536 -541 -528
rect -501 -536 -497 -528
rect -491 -536 -487 -528
rect -473 -536 -469 -528
rect -463 -536 -459 -528
rect -1169 -616 -1165 -608
rect -1157 -616 -1153 -608
rect -758 -612 -754 -604
rect -746 -612 -742 -604
rect -1222 -709 -1218 -701
rect -1212 -709 -1208 -701
rect -1194 -709 -1190 -701
rect -1184 -709 -1180 -701
rect -1139 -709 -1135 -701
rect -1129 -709 -1125 -701
rect -1111 -709 -1107 -701
rect -1101 -709 -1097 -701
rect -1032 -709 -1028 -701
rect -1022 -709 -1018 -701
rect -1004 -709 -1000 -701
rect -994 -709 -990 -701
rect -949 -709 -945 -701
rect -939 -709 -935 -701
rect -921 -709 -917 -701
rect -911 -709 -907 -701
<< m2contact >>
rect -1286 43 -1282 47
rect -819 43 -815 47
rect -855 38 -851 43
rect -1256 17 -1252 21
rect -1207 17 -1203 21
rect -1111 29 -1107 33
rect -1090 21 -1086 25
rect -1014 29 -1010 33
rect -936 29 -932 33
rect -864 21 -860 25
rect -1104 14 -1100 18
rect -441 38 -437 42
rect -700 29 -696 33
rect -680 22 -676 26
rect -604 29 -600 33
rect -1187 -1 -1183 3
rect -692 14 -688 18
rect -522 29 -518 33
rect -450 21 -446 25
rect -776 -1 -772 3
rect -1335 -9 -1331 -5
rect -1273 -19 -1269 -15
rect -1090 -16 -1086 -12
rect -1199 -26 -1195 -22
rect -1186 -34 -1182 -30
rect -680 -16 -676 -12
rect -788 -20 -784 -16
rect -775 -30 -771 -26
rect -1286 -149 -1282 -145
rect -819 -149 -815 -145
rect -855 -154 -851 -149
rect -1256 -175 -1252 -171
rect -1207 -175 -1203 -171
rect -1111 -163 -1107 -159
rect -1090 -171 -1086 -167
rect -1014 -163 -1010 -159
rect -936 -163 -932 -159
rect -864 -171 -860 -167
rect -1104 -178 -1100 -174
rect -441 -154 -437 -150
rect -700 -163 -696 -159
rect -680 -170 -676 -166
rect -604 -163 -600 -159
rect -1187 -193 -1183 -189
rect -692 -178 -688 -174
rect -522 -163 -518 -159
rect -450 -171 -446 -167
rect -776 -193 -772 -189
rect -1335 -201 -1331 -197
rect -1273 -211 -1269 -207
rect -1090 -208 -1086 -204
rect -1199 -218 -1195 -214
rect -1186 -226 -1182 -222
rect -680 -208 -676 -204
rect -788 -212 -784 -208
rect -775 -222 -771 -218
rect -1286 -340 -1282 -336
rect -819 -340 -815 -336
rect -855 -345 -851 -340
rect -1256 -366 -1252 -362
rect -1207 -366 -1203 -362
rect -1111 -354 -1107 -350
rect -1090 -362 -1086 -358
rect -1014 -354 -1010 -350
rect -936 -354 -932 -350
rect -864 -362 -860 -358
rect -1104 -369 -1100 -365
rect -441 -345 -437 -341
rect -700 -354 -696 -350
rect -680 -361 -676 -357
rect -604 -354 -600 -350
rect -1187 -384 -1183 -380
rect -692 -369 -688 -365
rect -522 -354 -518 -350
rect -450 -362 -446 -358
rect -776 -384 -772 -380
rect -1335 -392 -1331 -388
rect -1273 -402 -1269 -398
rect -1090 -399 -1086 -395
rect -1199 -409 -1195 -405
rect -1186 -417 -1182 -413
rect -680 -399 -676 -395
rect -788 -403 -784 -399
rect -775 -413 -771 -409
rect -1287 -526 -1283 -522
rect -820 -526 -816 -522
rect -856 -531 -852 -526
rect -1257 -552 -1253 -548
rect -1208 -552 -1204 -548
rect -1112 -540 -1108 -536
rect -1091 -548 -1087 -544
rect -1015 -540 -1011 -536
rect -937 -540 -933 -536
rect -865 -548 -861 -544
rect -1105 -555 -1101 -551
rect -442 -531 -438 -527
rect -701 -540 -697 -536
rect -681 -547 -677 -543
rect -605 -540 -601 -536
rect -1188 -570 -1184 -566
rect -693 -555 -689 -551
rect -523 -540 -519 -536
rect -451 -548 -447 -544
rect -777 -570 -773 -566
rect -1335 -578 -1331 -574
rect -1274 -588 -1269 -584
rect -1297 -652 -1293 -648
rect -1091 -585 -1087 -581
rect -1200 -595 -1196 -591
rect -1187 -603 -1183 -599
rect -681 -585 -677 -581
rect -789 -589 -785 -585
rect -776 -599 -772 -595
rect -1053 -663 -1049 -659
rect -965 -703 -961 -699
rect -1239 -721 -1235 -717
rect -1152 -721 -1148 -717
rect -1297 -728 -1293 -724
rect -1086 -721 -1082 -717
rect -1053 -721 -1049 -717
rect -1073 -728 -1069 -724
rect -346 -667 -342 -663
rect -959 -741 -955 -737
rect -1335 -751 -1331 -747
<< psubstratepcontact >>
rect -1238 -3 -1234 1
rect -1132 -2 -1128 2
rect -1035 -3 -1031 1
rect -949 -2 -945 2
rect -875 -3 -871 1
rect -721 -3 -717 1
rect -625 -2 -621 2
rect -543 -2 -539 2
rect -461 -2 -457 2
rect -757 -77 -753 -73
rect -1168 -81 -1164 -77
rect -1238 -195 -1234 -191
rect -1132 -194 -1128 -190
rect -1035 -195 -1031 -191
rect -949 -194 -945 -190
rect -875 -195 -871 -191
rect -721 -195 -717 -191
rect -625 -194 -621 -190
rect -543 -194 -539 -190
rect -461 -194 -457 -190
rect -757 -269 -753 -265
rect -1168 -273 -1164 -269
rect -1238 -386 -1234 -382
rect -1132 -385 -1128 -381
rect -1035 -386 -1031 -382
rect -949 -385 -945 -381
rect -875 -386 -871 -382
rect -721 -386 -717 -382
rect -625 -385 -621 -381
rect -543 -385 -539 -381
rect -461 -385 -457 -381
rect -757 -460 -753 -456
rect -1168 -464 -1164 -460
rect -1239 -572 -1235 -568
rect -1133 -571 -1129 -567
rect -1036 -572 -1032 -568
rect -950 -571 -946 -567
rect -876 -572 -872 -568
rect -722 -572 -718 -568
rect -626 -571 -622 -567
rect -544 -571 -540 -567
rect -462 -571 -458 -567
rect -758 -646 -754 -642
rect -1169 -650 -1165 -646
rect -1183 -745 -1179 -741
rect -1100 -745 -1096 -741
rect -993 -745 -989 -741
rect -910 -745 -906 -741
<< nsubstratencontact >>
rect -1238 44 -1234 48
rect -1223 44 -1219 48
rect -1171 45 -1167 49
rect -1163 45 -1159 49
rect -1153 45 -1149 49
rect -1143 45 -1139 49
rect -1133 45 -1129 49
rect -1074 45 -1070 49
rect -1066 45 -1062 49
rect -1056 45 -1052 49
rect -1046 45 -1042 49
rect -1036 45 -1032 49
rect -988 45 -984 49
rect -980 45 -976 49
rect -970 45 -966 49
rect -960 45 -956 49
rect -950 45 -946 49
rect -914 45 -910 49
rect -906 45 -902 49
rect -896 45 -892 49
rect -886 45 -882 49
rect -876 45 -872 49
rect -760 45 -756 49
rect -752 45 -748 49
rect -742 45 -738 49
rect -732 45 -728 49
rect -722 45 -718 49
rect -664 45 -660 49
rect -656 45 -652 49
rect -646 45 -642 49
rect -636 45 -632 49
rect -626 45 -622 49
rect -582 45 -578 49
rect -574 45 -570 49
rect -564 45 -560 49
rect -554 45 -550 49
rect -544 45 -540 49
rect -500 45 -496 49
rect -492 45 -488 49
rect -482 45 -478 49
rect -472 45 -468 49
rect -462 45 -458 49
rect -757 -30 -753 -26
rect -742 -30 -738 -26
rect -1168 -34 -1164 -30
rect -1153 -34 -1149 -30
rect -1238 -148 -1234 -144
rect -1223 -148 -1219 -144
rect -1171 -147 -1167 -143
rect -1163 -147 -1159 -143
rect -1153 -147 -1149 -143
rect -1143 -147 -1139 -143
rect -1133 -147 -1129 -143
rect -1074 -147 -1070 -143
rect -1066 -147 -1062 -143
rect -1056 -147 -1052 -143
rect -1046 -147 -1042 -143
rect -1036 -147 -1032 -143
rect -988 -147 -984 -143
rect -980 -147 -976 -143
rect -970 -147 -966 -143
rect -960 -147 -956 -143
rect -950 -147 -946 -143
rect -914 -147 -910 -143
rect -906 -147 -902 -143
rect -896 -147 -892 -143
rect -886 -147 -882 -143
rect -876 -147 -872 -143
rect -760 -147 -756 -143
rect -752 -147 -748 -143
rect -742 -147 -738 -143
rect -732 -147 -728 -143
rect -722 -147 -718 -143
rect -664 -147 -660 -143
rect -656 -147 -652 -143
rect -646 -147 -642 -143
rect -636 -147 -632 -143
rect -626 -147 -622 -143
rect -582 -147 -578 -143
rect -574 -147 -570 -143
rect -564 -147 -560 -143
rect -554 -147 -550 -143
rect -544 -147 -540 -143
rect -500 -147 -496 -143
rect -492 -147 -488 -143
rect -482 -147 -478 -143
rect -472 -147 -468 -143
rect -462 -147 -458 -143
rect -757 -222 -753 -218
rect -742 -222 -738 -218
rect -1168 -226 -1164 -222
rect -1153 -226 -1149 -222
rect -1238 -339 -1234 -335
rect -1223 -339 -1219 -335
rect -1171 -338 -1167 -334
rect -1163 -338 -1159 -334
rect -1153 -338 -1149 -334
rect -1143 -338 -1139 -334
rect -1133 -338 -1129 -334
rect -1074 -338 -1070 -334
rect -1066 -338 -1062 -334
rect -1056 -338 -1052 -334
rect -1046 -338 -1042 -334
rect -1036 -338 -1032 -334
rect -988 -338 -984 -334
rect -980 -338 -976 -334
rect -970 -338 -966 -334
rect -960 -338 -956 -334
rect -950 -338 -946 -334
rect -914 -338 -910 -334
rect -906 -338 -902 -334
rect -896 -338 -892 -334
rect -886 -338 -882 -334
rect -876 -338 -872 -334
rect -760 -338 -756 -334
rect -752 -338 -748 -334
rect -742 -338 -738 -334
rect -732 -338 -728 -334
rect -722 -338 -718 -334
rect -664 -338 -660 -334
rect -656 -338 -652 -334
rect -646 -338 -642 -334
rect -636 -338 -632 -334
rect -626 -338 -622 -334
rect -582 -338 -578 -334
rect -574 -338 -570 -334
rect -564 -338 -560 -334
rect -554 -338 -550 -334
rect -544 -338 -540 -334
rect -500 -338 -496 -334
rect -492 -338 -488 -334
rect -482 -338 -478 -334
rect -472 -338 -468 -334
rect -462 -338 -458 -334
rect -757 -413 -753 -409
rect -742 -413 -738 -409
rect -1168 -417 -1164 -413
rect -1153 -417 -1149 -413
rect -1239 -525 -1235 -521
rect -1224 -525 -1220 -521
rect -1172 -524 -1168 -520
rect -1164 -524 -1160 -520
rect -1154 -524 -1150 -520
rect -1144 -524 -1140 -520
rect -1134 -524 -1130 -520
rect -1075 -524 -1071 -520
rect -1067 -524 -1063 -520
rect -1057 -524 -1053 -520
rect -1047 -524 -1043 -520
rect -1037 -524 -1033 -520
rect -989 -524 -985 -520
rect -981 -524 -977 -520
rect -971 -524 -967 -520
rect -961 -524 -957 -520
rect -951 -524 -947 -520
rect -915 -524 -911 -520
rect -907 -524 -903 -520
rect -897 -524 -893 -520
rect -887 -524 -883 -520
rect -877 -524 -873 -520
rect -761 -524 -757 -520
rect -753 -524 -749 -520
rect -743 -524 -739 -520
rect -733 -524 -729 -520
rect -723 -524 -719 -520
rect -665 -524 -661 -520
rect -657 -524 -653 -520
rect -647 -524 -643 -520
rect -637 -524 -633 -520
rect -627 -524 -623 -520
rect -583 -524 -579 -520
rect -575 -524 -571 -520
rect -565 -524 -561 -520
rect -555 -524 -551 -520
rect -545 -524 -541 -520
rect -501 -524 -497 -520
rect -493 -524 -489 -520
rect -483 -524 -479 -520
rect -473 -524 -469 -520
rect -463 -524 -459 -520
rect -758 -599 -754 -595
rect -743 -599 -739 -595
rect -1169 -603 -1165 -599
rect -1154 -603 -1150 -599
rect -1222 -697 -1218 -693
rect -1214 -697 -1210 -693
rect -1204 -697 -1200 -693
rect -1194 -697 -1190 -693
rect -1184 -697 -1180 -693
rect -1139 -697 -1135 -693
rect -1131 -697 -1127 -693
rect -1121 -697 -1117 -693
rect -1111 -697 -1107 -693
rect -1101 -697 -1097 -693
rect -1032 -697 -1028 -693
rect -1024 -697 -1020 -693
rect -1014 -697 -1010 -693
rect -1004 -697 -1000 -693
rect -994 -697 -990 -693
rect -949 -697 -945 -693
rect -941 -697 -937 -693
rect -931 -697 -927 -693
rect -921 -697 -917 -693
rect -911 -697 -907 -693
<< labels >>
rlabel pdcontact -461 -530 -461 -530 1 M7source
rlabel pdcontact -501 -529 -501 -529 1 M6source
rlabel pdcontact -543 -530 -543 -530 1 M7source
rlabel pdcontact -583 -529 -583 -529 1 M6source
rlabel pdcontact -625 -530 -625 -530 1 M7source
rlabel pdcontact -665 -529 -665 -529 1 M6source
rlabel pdcontact -721 -530 -721 -530 1 M7source
rlabel pdcontact -761 -529 -761 -529 1 M6source
rlabel pdcontact -875 -530 -875 -530 1 M7source
rlabel pdcontact -915 -529 -915 -529 1 M6source
rlabel pdcontact -949 -530 -949 -530 1 M7source
rlabel pdcontact -989 -529 -989 -529 1 M6source
rlabel pdcontact -1035 -530 -1035 -530 1 M7source
rlabel pdcontact -1075 -529 -1075 -529 1 M6source
rlabel pdcontact -1132 -530 -1132 -530 1 M7source
rlabel pdcontact -1172 -529 -1172 -529 1 M6source
rlabel metal1 -1356 -510 -1356 -506 3 vdd!
rlabel metal1 -384 -561 -384 -557 7 FF1
rlabel metal2 -1320 -607 -1316 -607 1 clock
rlabel metal2 -1335 -806 -1331 -806 1 gnd!
rlabel metal1 -1297 -590 -1293 -590 1 D
rlabel pdcontact -1099 -703 -1099 -703 1 M7source
rlabel pdcontact -1139 -702 -1139 -702 1 M6source
rlabel pdcontact -1182 -703 -1182 -703 1 M7source
rlabel pdcontact -1222 -702 -1222 -702 1 M6source
rlabel pdcontact -909 -703 -909 -703 1 M7source
rlabel pdcontact -949 -702 -949 -702 1 M6source
rlabel pdcontact -992 -703 -992 -703 1 M7source
rlabel pdcontact -1032 -702 -1032 -702 1 M6source
rlabel pdcontact -460 -344 -460 -344 1 M7source
rlabel pdcontact -500 -343 -500 -343 1 M6source
rlabel pdcontact -542 -344 -542 -344 1 M7source
rlabel pdcontact -582 -343 -582 -343 1 M6source
rlabel pdcontact -624 -344 -624 -344 1 M7source
rlabel pdcontact -664 -343 -664 -343 1 M6source
rlabel pdcontact -720 -344 -720 -344 1 M7source
rlabel pdcontact -760 -343 -760 -343 1 M6source
rlabel pdcontact -874 -344 -874 -344 1 M7source
rlabel pdcontact -914 -343 -914 -343 1 M6source
rlabel pdcontact -948 -344 -948 -344 1 M7source
rlabel pdcontact -988 -343 -988 -343 1 M6source
rlabel pdcontact -1034 -344 -1034 -344 1 M7source
rlabel pdcontact -1074 -343 -1074 -343 1 M6source
rlabel pdcontact -1131 -344 -1131 -344 1 M7source
rlabel pdcontact -1171 -343 -1171 -343 1 M6source
rlabel metal1 -385 -375 -385 -371 1 FF2
rlabel pdcontact -460 -153 -460 -153 1 M7source
rlabel pdcontact -500 -152 -500 -152 1 M6source
rlabel pdcontact -542 -153 -542 -153 1 M7source
rlabel pdcontact -582 -152 -582 -152 1 M6source
rlabel pdcontact -624 -153 -624 -153 1 M7source
rlabel pdcontact -664 -152 -664 -152 1 M6source
rlabel pdcontact -720 -153 -720 -153 1 M7source
rlabel pdcontact -760 -152 -760 -152 1 M6source
rlabel pdcontact -874 -153 -874 -153 1 M7source
rlabel pdcontact -914 -152 -914 -152 1 M6source
rlabel pdcontact -948 -153 -948 -153 1 M7source
rlabel pdcontact -988 -152 -988 -152 1 M6source
rlabel pdcontact -1034 -153 -1034 -153 1 M7source
rlabel pdcontact -1074 -152 -1074 -152 1 M6source
rlabel pdcontact -1131 -153 -1131 -153 1 M7source
rlabel pdcontact -1171 -152 -1171 -152 1 M6source
rlabel metal1 -385 -184 -385 -180 1 FF3
rlabel pdcontact -460 39 -460 39 1 M7source
rlabel pdcontact -500 40 -500 40 1 M6source
rlabel pdcontact -542 39 -542 39 1 M7source
rlabel pdcontact -582 40 -582 40 1 M6source
rlabel pdcontact -624 39 -624 39 1 M7source
rlabel pdcontact -664 40 -664 40 1 M6source
rlabel pdcontact -720 39 -720 39 1 M7source
rlabel pdcontact -760 40 -760 40 1 M6source
rlabel pdcontact -874 39 -874 39 1 M7source
rlabel pdcontact -914 40 -914 40 1 M6source
rlabel pdcontact -948 39 -948 39 1 M7source
rlabel pdcontact -988 40 -988 40 1 M6source
rlabel pdcontact -1034 39 -1034 39 1 M7source
rlabel pdcontact -1074 40 -1074 40 1 M6source
rlabel pdcontact -1131 39 -1131 39 1 M7source
rlabel pdcontact -1171 40 -1171 40 1 M6source
rlabel metal1 -413 8 -413 12 1 FF4
<< end >>
