spice test
M1000 out vin vdd vdd pfet w=7 l=2
+ ad=49 pd=28 as=49 ps=28
M1001 out vin gnd gnd nfet w=4 l=2
+ ad=32 pd=24 as=32 ps=24
vdd vdd gnd 5
vin vin gnd 5
rgnd gnd 0 1e-6
.model nfet NMOS LEVEL=3 PHI=0.600000 TOX=2.1200E-08
+ XJ=0.200000U TPG=1 VTO=0.7860 DELTA=6.9670E-01
+ LD=1.6470E-07 KP=9.6379E-05 UO=591.7 THETA=8.1220E-02
+ RSH=8.5450E+01 GAMMA=0.5863 NSUB=1.6160E+16
+ NFS=5.0000E+12 VMAX=2.0820E+05 ETA=7.0660E-02
+ KAPPA=1.3960E-01 CGDO=4.0241E-10 CGSO=4.0241E-10
+ CGBO=3.6144E-10 CJ=3.8541E-04 MJ=1.1854
+ CJSW=1.3940E-10 MJSW=0.125195 PB=0.800000
.model pfet PMOS LEVEL=3 PHI=0.600000 TOX=2.1200E-08
+ XJ=0.200000U TPG=-1 VTO=-0.9056 DELTA=1.5200E+00
+ LD=2.2000E-08 KP=2.9352E-05 UO=180.2 THETA=1.2480E-01
+ RSH=1.0470E+02 GAMMA=0.4863 NSUB=1.8900E+16
+ NFS=3.46E+12 VMAX=3.7320E+05 ETA=1.6410E-01
+ KAPPA=9.6940E+00 CGDO=5.3752E-11 CGSO=5.3752E-11
+ CGBO=3.3650E-10 CJ=4.8447E-04 MJ=0.5027
+ CJSW=1.6457E-10 MJSW=0.217168 PB=0.850000
.print dc v(out)
.print dc vin
.trans 1ns 100ns
.end

