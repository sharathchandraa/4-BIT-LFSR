spice file for OR gate using NAND gates
M1000 a_n821_n13# A vdd vdd pfet w=8 l=2
+ ad=96 pd=56 as=288 ps=168
M1001 vdd A a_n821_n13# vdd pfet w=8 l=2
+ ad=0 pd=0 as=0 ps=0
M1002 out a_n821_n13# vdd vdd pfet w=8 l=2
+ ad=96 pd=56 as=0 ps=0
M1003 vdd a_n695_n14# out vdd pfet w=8 l=2
+ ad=0 pd=0 as=0 ps=0
M1004 a_n695_n14# B vdd vdd pfet w=8 l=2
+ ad=96 pd=56 as=0 ps=0
M1005 vdd B a_n695_n14# vdd pfet w=8 l=2
+ ad=0 pd=0 as=0 ps=0
M1006 a_n812_n12# A a_n821_n13# Gnd nfet w=4 l=2
+ ad=64 pd=48 as=32 ps=24
M1007 gnd A a_n812_n12# Gnd nfet w=4 l=2
+ ad=96 pd=72 as=0 ps=0
M1008 a_n721_n12# a_n821_n13# out Gnd nfet w=4 l=2
+ ad=64 pd=48 as=32 ps=24
M1009 gnd a_n695_n14# a_n721_n12# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0
M1010 a_n639_n12# B a_n695_n14# Gnd nfet w=4 l=2
+ ad=64 pd=48 as=32 ps=24
M1011 gnd B a_n639_n12# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0
rgnd gnd 0 1e-6
v3 vdd gnd 5
v1 A 0 pulse(0 5 90ns 0ns 0ns 20ns 100ns)
v2 B 0 pulse(0 5 90ns 0ns 0ns 20ns 100ns)

.trans 1ns 300ns
..MODEL nfet NMOS ( kp=4.32e-4 vt0=0.4)
.MODEL pfet pMOS ( kp=1.12e-4 vt0=-0.4)

.print dc v(A)
.print dc v(B)
.print dc v(out)
.end

