* SPICE3 file created from OR.ext - technology: scmos

.option scale=1u

M1000 a_n821_n13# A vdd vdd pfet w=8 l=2
+ ad=96 pd=56 as=288 ps=168
M1001 vdd A a_n821_n13# vdd pfet w=8 l=2
+ ad=0 pd=0 as=0 ps=0
M1002 out a_n821_n13# vdd vdd pfet w=8 l=2
+ ad=96 pd=56 as=0 ps=0
M1003 vdd a_n695_n14# out vdd pfet w=8 l=2
+ ad=0 pd=0 as=0 ps=0
M1004 a_n695_n14# B vdd vdd pfet w=8 l=2
+ ad=96 pd=56 as=0 ps=0
M1005 vdd B a_n695_n14# vdd pfet w=8 l=2
+ ad=0 pd=0 as=0 ps=0
M1006 a_n812_n12# A a_n821_n13# Gnd nfet w=4 l=2
+ ad=64 pd=48 as=32 ps=24
M1007 gnd A a_n812_n12# Gnd nfet w=4 l=2
+ ad=96 pd=72 as=0 ps=0
M1008 a_n721_n12# a_n821_n13# out Gnd nfet w=4 l=2
+ ad=64 pd=48 as=32 ps=24
M1009 gnd a_n695_n14# a_n721_n12# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0
M1010 a_n639_n12# B a_n695_n14# Gnd nfet w=4 l=2
+ ad=64 pd=48 as=32 ps=24
M1011 gnd B a_n639_n12# Gnd nfet w=4 l=2
+ ad=0 pd=0 as=0 ps=0

